module top_1
#( parameter param177 = (((({(8'h9e)} ? {(8'hbc), (8'haf)} : ((8'hb2) == (8'hb4))) | (((8'h9c) ? (8'hb1) : (8'hb3)) ~^ (^(8'ha1)))) < ({(&(8'ha9)), {(8'hb8)}} <= {(~(8'had))})) * ((~|(((8'hb4) - (8'hb3)) ? ((8'hba) < (8'hb8)) : ((8'hb3) && (8'hab)))) + (((&(8'haf)) ? (+(7'h42)) : ((8'ha8) ? (8'hae) : (8'hb8))) < (((8'hb9) >> (8'ha1)) ? (~(8'hbf)) : ((8'hab) ? (8'had) : (8'hb0))))))
, parameter param178 = (param177 & param177) )
(y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'he8):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire4;
  input wire [(4'hb):(1'h0)] wire3;
  input wire signed [(5'h13):(1'h0)] wire2;
  input wire [(5'h11):(1'h0)] wire1;
  input wire signed [(3'h7):(1'h0)] wire0;
  wire [(4'h8):(1'h0)] wire175;
  wire signed [(2'h3):(1'h0)] wire174;
  wire signed [(4'hf):(1'h0)] wire173;
  wire signed [(3'h4):(1'h0)] wire172;
  wire [(4'ha):(1'h0)] wire171;
  wire [(5'h15):(1'h0)] wire170;
  reg signed [(2'h3):(1'h0)] reg169 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg168 = (1'h0);
  reg [(3'h4):(1'h0)] reg167 = (1'h0);
  reg [(4'hd):(1'h0)] reg166 = (1'h0);
  reg [(4'h8):(1'h0)] reg165 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg164 = (1'h0);
  wire [(5'h15):(1'h0)] wire163;
  wire [(3'h4):(1'h0)] wire162;
  wire signed [(4'hb):(1'h0)] wire161;
  wire [(4'he):(1'h0)] wire159;
  wire [(4'hb):(1'h0)] wire26;
  wire signed [(5'h10):(1'h0)] wire7;
  wire signed [(4'hf):(1'h0)] wire6;
  wire [(5'h12):(1'h0)] wire5;
  assign y = {wire175,
                 wire174,
                 wire173,
                 wire172,
                 wire171,
                 wire170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 wire163,
                 wire162,
                 wire161,
                 wire159,
                 wire26,
                 wire7,
                 wire6,
                 wire5,
                 (1'h0)};
  assign wire5 = ((8'hb3) > ($unsigned((wire2 ?
                     wire1[(4'hb):(2'h3)] : wire0[(1'h1):(1'h0)])) ^~ ((|$unsigned(wire3)) | (8'hb6))));
  assign wire6 = (($signed($signed(wire2)) * (|wire4[(3'h6):(1'h0)])) + (~(-wire5)));
  assign wire7 = wire0;
  module8_1 modinst27 (wire26, clk, wire3, wire6, wire0, wire4);
  module28_1 modinst160 (.clk(clk), .wire32(wire1), .wire31(wire26), .wire30(wire6), .y(wire159), .wire29(wire5));
  assign wire161 = wire0;
  assign wire162 = wire7;
  assign wire163 = $signed((^{{(wire0 ? wire26 : wire2)},
                       $unsigned((wire5 ? wire162 : wire159))}));
  always
    @(posedge clk) begin
      if (wire3[(1'h1):(1'h0)])
        begin
          if ((+$signed(wire4[(2'h2):(2'h2)])))
            begin
              reg164 <= wire6[(4'hc):(2'h2)];
            end
          else
            begin
              reg164 <= ((8'hab) ?
                  $unsigned(wire159[(4'he):(1'h0)]) : $signed($unsigned(wire3[(4'ha):(3'h7)])));
              reg165 <= wire6[(2'h3):(2'h2)];
              reg166 <= $unsigned((~&(|$unsigned($signed(wire163)))));
            end
          reg167 <= ($signed((^(wire5 <<< (~&wire159)))) ?
              $signed((|(wire3[(2'h2):(1'h1)] ?
                  (wire162 ?
                      (8'hb3) : (8'hac)) : wire5))) : {(wire7 || (+(8'ha8))),
                  ($unsigned($unsigned(wire6)) << (~(wire4 < wire4)))});
          reg168 <= ({{$unsigned(((8'hbb) ? wire5 : wire163))},
              {$unsigned($signed(reg166))}} < ($signed(wire5) & $signed(reg164[(3'h4):(1'h0)])));
          reg169 <= $signed(wire161[(3'h6):(3'h6)]);
        end
      else
        begin
          reg164 <= wire159[(4'h8):(3'h4)];
          reg165 <= {$unsigned((wire26[(3'h5):(1'h1)] ^~ ($unsigned(wire4) ^~ wire6))),
              (~((8'ha7) != (wire5[(4'hf):(2'h2)] ?
                  (wire7 <<< (8'h9e)) : (-wire0))))};
          reg166 <= (wire161 ~^ $unsigned((8'hab)));
        end
    end
  assign wire170 = $unsigned((^(8'hb2)));
  assign wire171 = ($unsigned({wire159[(4'hc):(2'h3)],
                       $unsigned((~(8'hb2)))}) <<< ($unsigned($unsigned($signed(reg168))) ?
                       wire3[(1'h1):(1'h1)] : (8'hbb)));
  assign wire172 = ($unsigned((~reg167)) + wire4[(3'h4):(2'h2)]);
  assign wire173 = $signed((reg169[(1'h0):(1'h0)] >> (reg168[(1'h0):(1'h0)] << ((wire171 < wire26) + {wire170,
                       reg169}))));
  assign wire174 = (8'hab);
  module28_1 modinst176 (wire175, clk, reg166, wire159, wire26, wire4);
endmodule

module module28_1  (y, clk, wire29, wire30, wire31, wire32);
  output wire [(32'h150):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire29;
  input wire signed [(4'h8):(1'h0)] wire30;
  input wire signed [(4'hb):(1'h0)] wire31;
  input wire [(5'h11):(1'h0)] wire32;
  wire [(2'h2):(1'h0)] wire158;
  wire [(4'ha):(1'h0)] wire156;
  wire [(5'h14):(1'h0)] wire131;
  wire [(3'h5):(1'h0)] wire130;
  wire signed [(5'h14):(1'h0)] wire129;
  wire [(2'h2):(1'h0)] wire128;
  wire [(5'h13):(1'h0)] wire126;
  wire [(2'h2):(1'h0)] wire104;
  wire [(4'h9):(1'h0)] wire103;
  wire signed [(4'hc):(1'h0)] wire102;
  wire signed [(4'hd):(1'h0)] wire101;
  wire [(2'h2):(1'h0)] wire33;
  reg [(5'h11):(1'h0)] reg34 = (1'h0);
  reg [(5'h15):(1'h0)] reg35 = (1'h0);
  reg [(2'h3):(1'h0)] reg36 = (1'h0);
  reg [(5'h10):(1'h0)] reg37 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg38 = (1'h0);
  reg [(5'h15):(1'h0)] reg39 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg40 = (1'h0);
  reg [(5'h12):(1'h0)] reg41 = (1'h0);
  reg [(4'ha):(1'h0)] reg42 = (1'h0);
  reg [(5'h14):(1'h0)] reg43 = (1'h0);
  reg [(4'hf):(1'h0)] reg44 = (1'h0);
  reg [(5'h13):(1'h0)] reg45 = (1'h0);
  wire [(4'hc):(1'h0)] wire67;
  wire signed [(5'h15):(1'h0)] wire69;
  wire [(2'h3):(1'h0)] wire99;
  assign y = {wire158,
                 wire156,
                 wire131,
                 wire130,
                 wire129,
                 wire128,
                 wire126,
                 wire104,
                 wire103,
                 wire102,
                 wire101,
                 wire33,
                 reg34,
                 reg35,
                 reg36,
                 reg37,
                 reg38,
                 reg39,
                 reg40,
                 reg41,
                 reg42,
                 reg43,
                 reg44,
                 reg45,
                 wire67,
                 wire69,
                 wire99,
                 (1'h0)};
  assign wire33 = $unsigned((^((~&(~wire32)) * (~&(!wire29)))));
  always
    @(posedge clk) begin
      if ({{(8'ha0)}})
        begin
          if ({wire33[(1'h1):(1'h1)]})
            begin
              reg34 <= $signed($unsigned($unsigned((~|{wire30}))));
              reg35 <= $unsigned(wire31[(1'h1):(1'h1)]);
              reg36 <= $signed(wire32);
              reg37 <= $unsigned({((^((7'h44) ? reg34 : reg35)) ?
                      ((~^wire29) > wire33[(1'h0):(1'h0)]) : wire32[(4'hb):(2'h2)])});
            end
          else
            begin
              reg34 <= reg37;
              reg35 <= $signed(($unsigned(wire33) ?
                  ($unsigned((reg35 == wire30)) ?
                      wire31 : $unsigned((wire31 ?
                          (8'haf) : reg36))) : (wire31 ?
                      (reg35[(1'h1):(1'h0)] * (reg37 ?
                          wire31 : reg35)) : $unsigned((reg36 || reg37)))));
            end
        end
      else
        begin
          if ($unsigned((^~(reg34[(2'h3):(1'h1)] * (&wire31[(1'h1):(1'h1)])))))
            begin
              reg34 <= $signed(wire33[(2'h2):(2'h2)]);
              reg35 <= $unsigned((!(8'haf)));
            end
          else
            begin
              reg34 <= wire31;
              reg35 <= wire31;
              reg36 <= (wire32 ~^ {reg36, $unsigned($signed(reg35))});
              reg37 <= wire30;
            end
          reg38 <= (~^$unsigned($unsigned(wire33)));
          reg39 <= wire30;
          reg40 <= (wire33 >= (+((|(-reg39)) | (((8'h9f) ?
              reg37 : wire31) ~^ {reg37}))));
          reg41 <= (-wire31);
        end
      reg42 <= reg38;
      reg43 <= $unsigned($unsigned(($unsigned(wire30) ?
          (^~((7'h41) - reg35)) : (wire31[(3'h4):(3'h4)] ?
              (8'haa) : $unsigned(reg36)))));
      reg44 <= (+(~^{(wire33[(1'h0):(1'h0)] ?
              wire33[(2'h2):(2'h2)] : wire31[(3'h5):(3'h5)]),
          $unsigned($signed(reg43))}));
      reg45 <= (((&reg44) ? reg39 : reg36) != wire32);
    end
  module46_1 modinst68 (wire67, clk, wire31, reg42, wire30, reg38);
  assign wire69 = (((wire67[(1'h0):(1'h0)] ? reg37 : reg42[(3'h4):(3'h4)]) ?
                          $unsigned(reg41[(1'h0):(1'h0)]) : (8'hb3)) ?
                      wire30[(1'h0):(1'h0)] : ($signed({{wire67, (7'h42)},
                              reg45[(2'h3):(1'h1)]}) ?
                          (~&$unsigned({reg38})) : ($unsigned($signed(wire32)) ?
                              wire33 : wire33[(1'h1):(1'h0)])));
  module70_1 modinst100 (wire99, clk, wire29, reg41, wire69, reg35, reg38);
  assign wire101 = (~|$unsigned((^~wire69[(4'ha):(1'h0)])));
  assign wire102 = $unsigned(reg41);
  assign wire103 = $unsigned(reg44);
  assign wire104 = reg44[(4'h8):(2'h2)];
  module105_1 modinst127 (.wire108(wire102), .y(wire126), .clk(clk), .wire107(wire103), .wire109(reg38), .wire106(reg35));
  assign wire128 = $signed((8'hbc));
  assign wire129 = reg40[(3'h5):(2'h2)];
  assign wire130 = $unsigned($signed(($unsigned(((8'hb4) ? wire30 : wire101)) ?
                       (!$signed(wire30)) : $signed({wire33}))));
  assign wire131 = ($signed((($signed(wire99) ?
                           $unsigned(wire31) : $signed((8'ha8))) != wire67)) ?
                       {(+{(8'hb0)}),
                           $signed(((reg38 ? reg39 : wire32) ?
                               (~&reg37) : (~&wire32)))} : wire32[(3'h5):(1'h1)]);
  module132_1 modinst157 (.clk(clk), .wire134(reg44), .wire136(wire30), .wire135(wire69), .y(wire156), .wire133(reg39));
  assign wire158 = (((-(~&wire103[(4'h8):(4'h8)])) ?
                       wire126 : wire102) < reg41[(5'h11):(5'h11)]);
endmodule

module module8_1
#(parameter param25 = (8'hbd))
(y, clk, wire12, wire11, wire10, wire9);
  output wire [(32'h7c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h6):(1'h0)] wire12;
  input wire [(4'hf):(1'h0)] wire11;
  input wire [(3'h7):(1'h0)] wire10;
  input wire [(4'ha):(1'h0)] wire9;
  wire signed [(4'hd):(1'h0)] wire24;
  wire [(4'ha):(1'h0)] wire23;
  wire [(5'h15):(1'h0)] wire22;
  wire signed [(3'h4):(1'h0)] wire21;
  wire [(4'hd):(1'h0)] wire20;
  wire signed [(5'h14):(1'h0)] wire19;
  reg [(5'h10):(1'h0)] reg18 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg17 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire16;
  wire signed [(2'h3):(1'h0)] wire15;
  wire [(2'h2):(1'h0)] wire14;
  wire [(3'h6):(1'h0)] wire13;
  assign y = {wire24,
                 wire23,
                 wire22,
                 wire21,
                 wire20,
                 wire19,
                 reg18,
                 reg17,
                 wire16,
                 wire15,
                 wire14,
                 wire13,
                 (1'h0)};
  assign wire13 = (wire11 + $signed((((wire12 <<< wire10) ?
                      wire12 : $signed(wire11)) == (!(wire9 | (8'ha7))))));
  assign wire14 = (~$signed(((-wire12[(2'h2):(1'h0)]) + $unsigned((wire12 * wire12)))));
  assign wire15 = wire11;
  assign wire16 = wire11;
  always
    @(posedge clk) begin
      reg17 <= (wire14 << (wire16[(2'h3):(1'h1)] >> $signed($unsigned(((8'hba) < wire16)))));
      reg18 <= ($signed((&$unsigned($unsigned(wire15)))) ?
          $unsigned({wire11[(4'h8):(3'h4)]}) : wire16);
    end
  assign wire19 = ($unsigned({(7'h40)}) ?
                      $signed(wire16) : reg18[(4'ha):(4'h8)]);
  assign wire20 = {((wire11[(4'hc):(4'hb)] ~^ wire16) << $unsigned($unsigned(wire9))),
                      (($signed((!wire11)) ?
                          wire15 : wire13) ^~ {reg17[(2'h2):(2'h2)]})};
  assign wire21 = (~|(wire14 ?
                      $signed($unsigned((wire9 - wire15))) : reg17[(2'h3):(2'h2)]));
  assign wire22 = ({$unsigned((((8'ha4) ?
                          (7'h43) : wire19) >>> (!(8'ha4))))} < (wire14 | (~|$unsigned(wire11[(4'hd):(3'h7)]))));
  assign wire23 = (&$unsigned((|wire19)));
  assign wire24 = $unsigned(wire11[(3'h4):(1'h0)]);
endmodule

module module132_1  (y, clk, wire136, wire135, wire134, wire133);
  output wire [(32'hbf):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire136;
  input wire signed [(5'h15):(1'h0)] wire135;
  input wire [(4'h9):(1'h0)] wire134;
  input wire [(5'h13):(1'h0)] wire133;
  wire signed [(5'h10):(1'h0)] wire155;
  wire signed [(2'h2):(1'h0)] wire154;
  wire signed [(5'h12):(1'h0)] wire153;
  wire signed [(4'h9):(1'h0)] wire152;
  wire [(3'h6):(1'h0)] wire151;
  wire [(4'ha):(1'h0)] wire150;
  wire [(4'hb):(1'h0)] wire149;
  wire [(2'h3):(1'h0)] wire148;
  wire [(5'h11):(1'h0)] wire147;
  reg signed [(2'h2):(1'h0)] reg146 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg145 = (1'h0);
  reg [(5'h14):(1'h0)] reg144 = (1'h0);
  reg [(4'hc):(1'h0)] reg143 = (1'h0);
  reg [(2'h2):(1'h0)] reg142 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg141 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg140 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire139;
  wire signed [(4'h8):(1'h0)] wire138;
  wire signed [(4'he):(1'h0)] wire137;
  assign y = {wire155,
                 wire154,
                 wire153,
                 wire152,
                 wire151,
                 wire150,
                 wire149,
                 wire148,
                 wire147,
                 reg146,
                 reg145,
                 reg144,
                 reg143,
                 reg142,
                 reg141,
                 reg140,
                 wire139,
                 wire138,
                 wire137,
                 (1'h0)};
  assign wire137 = wire134;
  assign wire138 = ((|(~&(|wire137))) ?
                       wire135[(2'h2):(2'h2)] : ($unsigned((!$signed(wire133))) ?
                           (wire137[(4'he):(1'h1)] ?
                               {$unsigned(wire137)} : ($signed(wire135) * (wire136 <<< wire136))) : wire135));
  assign wire139 = {(-$signed(((wire135 ? wire133 : wire138) ?
                           $signed(wire135) : wire138[(4'h8):(4'h8)])))};
  always
    @(posedge clk) begin
      reg140 <= {$signed((~^wire137))};
      if (wire135)
        begin
          reg141 <= ((wire133 ? $unsigned((~^(+wire135))) : wire133) ?
              $unsigned({$unsigned((+wire137))}) : $unsigned((((+wire136) <= (&reg140)) ?
                  (^~(^wire139)) : $signed((wire134 ~^ wire136)))));
          reg142 <= reg140;
          reg143 <= $signed((~((wire133 ?
              (^~reg140) : $unsigned(wire134)) == (!wire134))));
        end
      else
        begin
          reg141 <= ($signed((7'h41)) ?
              {(($unsigned(reg141) ? $unsigned(wire139) : $signed(wire133)) ?
                      ($signed((8'ha4)) ~^ wire139) : (wire134 <= (+wire136)))} : ($signed(({wire135,
                  wire137} ^ reg141)) >= (~wire139[(4'h9):(4'h8)])));
        end
      reg144 <= $unsigned(($signed({wire137[(4'hb):(3'h6)],
          $unsigned(wire139)}) - (reg141 ?
          wire137 : {wire136[(3'h5):(2'h3)], {reg140, wire139}})));
      reg145 <= wire138[(2'h3):(1'h0)];
      reg146 <= ($unsigned({{reg144[(4'hd):(2'h2)],
              (~&reg141)}}) == (($signed({reg141}) != $signed(wire136[(3'h6):(3'h4)])) ?
          $signed(({wire134, (8'ha7)} && reg142[(2'h2):(2'h2)])) : (&reg141)));
    end
  assign wire147 = reg146[(2'h2):(2'h2)];
  assign wire148 = $signed(wire138);
  assign wire149 = ($unsigned($signed(wire136[(2'h3):(1'h1)])) ?
                       {((wire138[(2'h2):(2'h2)] ?
                               $signed(reg140) : reg144) != {$signed(reg143)}),
                           (($signed(wire148) ?
                               (wire148 ? wire133 : wire136) : {wire138,
                                   reg141}) + ((reg144 ^ wire136) ?
                               reg144[(4'hf):(4'h8)] : (wire139 || wire135)))} : $unsigned((wire137[(3'h7):(3'h7)] * {$signed(wire147),
                           (wire139 <<< (7'h41))})));
  assign wire150 = wire135[(3'h6):(1'h0)];
  assign wire151 = wire138;
  assign wire152 = ($unsigned($unsigned(((wire151 && wire136) ?
                           $unsigned((8'hbb)) : (~|reg143)))) ?
                       (reg140 != ($signed((wire135 >>> wire150)) && (~^$unsigned(reg145)))) : wire147[(4'he):(4'h9)]);
  assign wire153 = ((8'ha2) ?
                       ($unsigned($unsigned($signed(wire148))) >>> $unsigned((wire136[(2'h2):(2'h2)] > (+reg140)))) : $unsigned({(~^(reg141 ?
                               wire149 : wire152))}));
  assign wire154 = $signed($signed($signed($signed(wire133))));
  assign wire155 = {wire139[(1'h1):(1'h0)]};
endmodule

module module105_1
#( parameter param125 = (^(((8'hb3) ? ((~&(8'hb2)) || ((7'h40) ? (8'hbd) : (8'hbf))) : {((8'hbd) || (8'ha1))}) >= {(((8'h9f) == (8'ha2)) ? (~&(8'ha0)) : (~(8'hb4))), {((7'h43) & (8'h9d)), (~&(8'h9c))}})) )
(y, clk, wire109, wire108, wire107, wire106);
  output wire [(32'hb8):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire109;
  input wire [(3'h4):(1'h0)] wire108;
  input wire [(4'h9):(1'h0)] wire107;
  input wire signed [(4'he):(1'h0)] wire106;
  wire signed [(4'h8):(1'h0)] wire124;
  wire signed [(3'h6):(1'h0)] wire123;
  wire [(4'hf):(1'h0)] wire122;
  reg [(4'hc):(1'h0)] reg121 = (1'h0);
  reg [(4'hb):(1'h0)] reg120 = (1'h0);
  reg [(5'h14):(1'h0)] reg119 = (1'h0);
  reg [(4'hb):(1'h0)] reg118 = (1'h0);
  reg [(3'h6):(1'h0)] reg117 = (1'h0);
  reg [(4'hd):(1'h0)] reg116 = (1'h0);
  reg [(5'h13):(1'h0)] reg115 = (1'h0);
  reg [(5'h13):(1'h0)] reg114 = (1'h0);
  wire [(5'h11):(1'h0)] wire113;
  wire signed [(2'h3):(1'h0)] wire112;
  wire [(4'h9):(1'h0)] wire111;
  wire [(4'he):(1'h0)] wire110;
  assign y = {wire124,
                 wire123,
                 wire122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 reg117,
                 reg116,
                 reg115,
                 reg114,
                 wire113,
                 wire112,
                 wire111,
                 wire110,
                 (1'h0)};
  assign wire110 = $unsigned(($signed((~|$signed(wire106))) ?
                       wire107[(4'h8):(3'h6)] : wire108[(3'h4):(2'h3)]));
  assign wire111 = wire107;
  assign wire112 = $unsigned(((((wire108 ? wire106 : wire107) ?
                       (wire108 || wire108) : (~&wire108)) != ($unsigned(wire110) <<< wire109[(1'h0):(1'h0)])) << (+wire109[(4'hb):(2'h2)])));
  assign wire113 = $unsigned((~^({$signed(wire112)} ^ ((~&(8'hae)) ?
                       wire109[(4'h9):(1'h1)] : $signed((8'hbd))))));
  always
    @(posedge clk) begin
      if (((^(wire112 ?
              wire108 : ((&wire106) ? (~|wire111) : $signed(wire106)))) ?
          $unsigned(wire112[(2'h2):(1'h0)]) : $signed((wire110[(2'h2):(1'h0)] + (((8'h9c) & wire113) ^ {wire113,
              wire109})))))
        begin
          reg114 <= (~|((wire109 ? wire113 : $signed((|wire110))) ?
              {{wire108[(3'h4):(1'h1)]}, wire109} : (&(8'ha7))));
          reg115 <= $unsigned({($signed((wire112 ?
                  wire107 : wire107)) != wire109)});
          reg116 <= (((reg114 ?
                  (reg114[(4'hc):(1'h0)] ?
                      $signed((7'h44)) : $unsigned(wire111)) : {$unsigned(wire110)}) ~^ (^(7'h42))) ?
              $signed(reg115[(2'h2):(2'h2)]) : $signed(((8'hb0) ?
                  $unsigned(wire111[(4'h9):(2'h2)]) : wire113[(4'hd):(3'h6)])));
        end
      else
        begin
          reg114 <= $signed((!(~&$signed($signed(wire113)))));
          if (reg115[(5'h12):(5'h10)])
            begin
              reg115 <= wire106[(4'h8):(3'h6)];
              reg116 <= ($signed(wire113[(2'h3):(2'h2)]) * $signed($unsigned(((wire108 ?
                  reg116 : wire109) << (wire107 * wire108)))));
              reg117 <= ((^~{wire109[(4'hb):(3'h4)],
                  (~(wire110 == wire113))}) | $signed($signed($signed($signed(wire110)))));
              reg118 <= ((wire112[(2'h3):(1'h0)] << wire113[(1'h1):(1'h1)]) >> $signed(wire106));
            end
          else
            begin
              reg115 <= (~^((8'ha3) | $unsigned($signed((~&wire111)))));
              reg116 <= (wire108 >>> $unsigned(wire111));
              reg117 <= wire109[(1'h0):(1'h0)];
              reg118 <= reg116[(3'h5):(1'h0)];
            end
          reg119 <= $unsigned({wire109});
          reg120 <= ((+(({wire108, reg118} >>> (wire109 ?
                  reg117 : (8'hb3))) ~^ ((~^reg119) <= (reg119 ?
                  reg115 : wire107)))) ?
              $unsigned((wire108[(3'h4):(2'h3)] <= (^$unsigned(wire109)))) : {$unsigned({(8'hb6)}),
                  {reg118, (~|wire111[(2'h2):(1'h0)])}});
          reg121 <= wire108[(3'h4):(2'h2)];
        end
    end
  assign wire122 = $signed((reg121[(4'h9):(3'h7)] ?
                       reg120[(2'h3):(1'h0)] : {$unsigned((8'ha5)),
                           reg119[(4'hc):(3'h5)]}));
  assign wire123 = {$signed({reg116}),
                       ($unsigned($signed($unsigned(wire106))) <<< (8'ha8))};
  assign wire124 = (^~(^(8'hbd)));
endmodule

module module70_1  (y, clk, wire75, wire74, wire73, wire72, wire71);
  output wire [(32'hcc):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hc):(1'h0)] wire75;
  input wire [(5'h12):(1'h0)] wire74;
  input wire signed [(4'hd):(1'h0)] wire73;
  input wire [(2'h2):(1'h0)] wire72;
  input wire signed [(4'h8):(1'h0)] wire71;
  reg signed [(3'h4):(1'h0)] reg98 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg97 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire96;
  wire [(3'h6):(1'h0)] wire95;
  wire signed [(5'h12):(1'h0)] wire94;
  wire [(3'h5):(1'h0)] wire93;
  reg signed [(4'ha):(1'h0)] reg92 = (1'h0);
  reg [(4'hd):(1'h0)] reg91 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire90;
  wire signed [(3'h5):(1'h0)] wire89;
  wire [(3'h7):(1'h0)] wire88;
  wire [(2'h3):(1'h0)] wire87;
  wire signed [(3'h4):(1'h0)] wire86;
  reg [(4'he):(1'h0)] reg85 = (1'h0);
  reg [(4'h8):(1'h0)] reg84 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg83 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg82 = (1'h0);
  reg [(4'h8):(1'h0)] reg81 = (1'h0);
  reg [(3'h5):(1'h0)] reg80 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg79 = (1'h0);
  reg [(4'ha):(1'h0)] reg78 = (1'h0);
  reg [(4'hb):(1'h0)] reg77 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg76 = (1'h0);
  assign y = {reg98,
                 reg97,
                 wire96,
                 wire95,
                 wire94,
                 wire93,
                 reg92,
                 reg91,
                 wire90,
                 wire89,
                 wire88,
                 wire87,
                 wire86,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 reg80,
                 reg79,
                 reg78,
                 reg77,
                 reg76,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg76 <= (|(~$unsigned(((wire75 != wire71) && (wire71 ~^ (8'ha0))))));
      reg77 <= wire72[(1'h0):(1'h0)];
      reg78 <= (~^(&(8'hbf)));
    end
  always
    @(posedge clk) begin
      reg79 <= $signed((reg76[(3'h6):(1'h1)] < {$signed({wire74})}));
      reg80 <= ($signed($unsigned(reg76[(2'h2):(1'h1)])) ?
          wire73[(4'hc):(4'ha)] : ((($unsigned(reg79) ?
                  (8'hb8) : $unsigned(wire71)) ?
              $signed((wire74 >= reg76)) : wire73) != (((wire71 ?
              wire73 : reg77) <= (wire71 ^ wire71)) & wire73)));
      reg81 <= ($unsigned($unsigned(($signed(wire73) > ((8'hb9) & wire74)))) ?
          ((~|({wire73} << (^~wire72))) | ($unsigned(reg80) ?
              (reg77 + wire74[(4'h9):(2'h3)]) : ($unsigned((8'hb9)) > {reg78,
                  wire75}))) : $signed(($signed(wire72[(1'h1):(1'h1)]) <= ($unsigned((8'hb4)) ~^ (reg79 * wire73)))));
      if ((&$unsigned((reg81 ? ((^reg80) ? reg81 : {reg81}) : wire75))))
        begin
          reg82 <= (~&$unsigned(((|{(8'ha0)}) >>> $signed(wire73))));
          reg83 <= $signed(reg78[(2'h3):(1'h1)]);
        end
      else
        begin
          if (reg80)
            begin
              reg82 <= {reg78[(4'ha):(1'h1)],
                  ({wire75,
                      ($signed((8'hbf)) | (~|reg78))} & (reg83[(2'h2):(2'h2)] ?
                      (^(+wire72)) : (|(^~wire73))))};
              reg83 <= (-$unsigned((((wire72 ? reg81 : wire71) ?
                  reg79[(3'h5):(1'h1)] : $signed((8'ha9))) < $signed((^reg76)))));
              reg84 <= {{$unsigned((+wire72[(1'h0):(1'h0)])),
                      reg79[(4'h9):(3'h6)]}};
            end
          else
            begin
              reg82 <= $unsigned((!$unsigned((8'hb2))));
              reg83 <= $unsigned($unsigned(reg83[(3'h6):(2'h2)]));
              reg84 <= $unsigned($signed(wire73));
              reg85 <= $unsigned((~wire71[(1'h0):(1'h0)]));
            end
        end
    end
  assign wire86 = $unsigned(((8'ha0) ? wire74 : reg84));
  assign wire87 = ((~|{((8'ha0) ?
                          reg83 : reg84)}) ^~ (reg85[(3'h5):(2'h2)] != reg80));
  assign wire88 = reg83;
  assign wire89 = {(|wire87[(1'h1):(1'h1)]),
                      (reg85[(2'h2):(1'h0)] ?
                          reg84[(3'h5):(2'h2)] : {{(~reg84),
                                  (wire88 * reg78)}})};
  assign wire90 = {(8'ha9)};
  always
    @(posedge clk) begin
      reg91 <= (^~{$signed(wire74[(3'h6):(2'h2)])});
    end
  always
    @(posedge clk) begin
      reg92 <= ((($unsigned((!reg81)) > $unsigned(reg82[(2'h2):(1'h1)])) ?
          wire74 : wire74) & $unsigned($unsigned(reg81)));
    end
  assign wire93 = {reg79[(4'hd):(3'h5)],
                      ($signed(reg80[(1'h1):(1'h1)]) ?
                          wire88[(3'h7):(1'h0)] : (reg85[(1'h1):(1'h1)] ?
                              wire74[(3'h6):(1'h1)] : (^~wire73)))};
  assign wire94 = reg76;
  assign wire95 = $unsigned(reg92);
  assign wire96 = {$unsigned((wire74[(4'hd):(3'h6)] <<< (~^$unsigned(reg82)))),
                      ($unsigned((!{reg79,
                          (8'hb5)})) <<< ({$signed(wire72)} >>> ({reg76} ?
                          $unsigned(wire71) : (wire71 ? (8'h9d) : reg82))))};
  always
    @(posedge clk) begin
      reg97 <= ($unsigned(($signed({wire71}) << $unsigned((reg78 & reg80)))) >>> (|($signed((wire88 != reg77)) > $unsigned($unsigned(reg78)))));
      reg98 <= wire95;
    end
endmodule

module module46_1
#( parameter param66 = {{{((8'haa) >>> (~&(8'hac)))}, (~&((&(8'had)) | ((8'haf) != (8'ha4))))}, ((~{((8'ha7) ? (8'ha4) : (8'hb0)), (~&(8'ha5))}) || ((((8'hb1) ? (8'haf) : (8'hb8)) ? ((8'hb3) < (8'hac)) : ((8'hbc) ? (7'h41) : (8'hb3))) ? (8'hb1) : ((~|(8'ha7)) >>> ((8'hbc) || (8'hb4)))))} )
(y, clk, wire50, wire49, wire48, wire47);
  output wire [(32'hc3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hb):(1'h0)] wire50;
  input wire [(4'ha):(1'h0)] wire49;
  input wire [(3'h4):(1'h0)] wire48;
  input wire signed [(3'h4):(1'h0)] wire47;
  wire [(4'hc):(1'h0)] wire65;
  wire signed [(2'h3):(1'h0)] wire64;
  wire [(4'hd):(1'h0)] wire63;
  wire [(5'h11):(1'h0)] wire62;
  wire signed [(4'hf):(1'h0)] wire61;
  wire signed [(5'h11):(1'h0)] wire60;
  wire [(4'he):(1'h0)] wire59;
  wire [(4'h9):(1'h0)] wire58;
  wire signed [(5'h12):(1'h0)] wire57;
  reg signed [(4'he):(1'h0)] reg56 = (1'h0);
  wire [(4'h9):(1'h0)] wire55;
  wire [(4'he):(1'h0)] wire54;
  wire signed [(4'h9):(1'h0)] wire53;
  wire [(4'hc):(1'h0)] wire52;
  wire signed [(5'h12):(1'h0)] wire51;
  assign y = {wire65,
                 wire64,
                 wire63,
                 wire62,
                 wire61,
                 wire60,
                 wire59,
                 wire58,
                 wire57,
                 reg56,
                 wire55,
                 wire54,
                 wire53,
                 wire52,
                 wire51,
                 (1'h0)};
  assign wire51 = wire47[(1'h1):(1'h0)];
  assign wire52 = $signed($signed(((&$unsigned(wire51)) >> (7'h44))));
  assign wire53 = wire52[(3'h7):(3'h6)];
  assign wire54 = (+$unsigned(($signed(((8'hae) | wire52)) <<< ((|wire50) ~^ $signed((8'haa))))));
  assign wire55 = ($signed(wire54[(4'hc):(3'h5)]) ?
                      $signed((((^(8'hb5)) ?
                          $signed(wire48) : $unsigned(wire48)) >>> (((8'hb4) ?
                              wire50 : wire52) ?
                          $unsigned(wire49) : (wire53 <= wire49)))) : wire48[(3'h4):(2'h2)]);
  always
    @(posedge clk) begin
      reg56 <= (wire52 && $unsigned((|((|wire53) ?
          {wire50} : (wire52 == wire47)))));
    end
  assign wire57 = (wire54 == $signed((|reg56)));
  assign wire58 = ($signed(wire55) ?
                      $signed({wire55, wire51}) : $unsigned(reg56));
  assign wire59 = reg56;
  assign wire60 = $unsigned((wire48[(1'h1):(1'h0)] ?
                      wire54[(4'hd):(3'h7)] : ((&(~|wire58)) << wire59)));
  assign wire61 = (wire55[(1'h1):(1'h0)] + (&{(~&(wire58 ? reg56 : wire52))}));
  assign wire62 = (wire50[(3'h6):(3'h6)] ?
                      $unsigned($signed(((~^wire49) ?
                          wire57[(4'hd):(4'hd)] : wire52[(2'h2):(2'h2)]))) : (wire49[(1'h0):(1'h0)] + (($unsigned(wire49) - (~^wire53)) | ((wire52 < wire50) ?
                          $signed(reg56) : wire47[(1'h1):(1'h1)]))));
  assign wire63 = wire51;
  assign wire64 = wire51;
  assign wire65 = ($unsigned((({wire54} ?
                          $signed(wire59) : wire54) >> (+$signed((8'ha6))))) ?
                      $signed((-($signed(wire64) ?
                          $signed(wire52) : wire47[(2'h3):(1'h0)]))) : wire50);
endmodule