module top
#( parameter param227 = (!(((^((8'ha7) ? (8'ha2) : (7'h41))) ? (((8'haf) ? (8'hb1) : (8'h9e)) >>> (&(7'h40))) : (((8'hbe) ? (7'h42) : (8'hb6)) ? {(8'hb6)} : {(8'h9f), (8'hb5)})) & (|(!(!(8'ha7)))))) )
(y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h21c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire3;
  input wire signed [(5'h14):(1'h0)] wire2;
  input wire signed [(4'hc):(1'h0)] wire1;
  input wire [(5'h13):(1'h0)] wire0;
  reg [(4'ha):(1'h0)] reg226 = (1'h0);
  reg [(4'hd):(1'h0)] reg225 = (1'h0);
  reg [(5'h12):(1'h0)] reg224 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg223 = (1'h0);
  reg [(4'h9):(1'h0)] reg222 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg221 = (1'h0);
  reg [(3'h7):(1'h0)] reg220 = (1'h0);
  wire [(3'h7):(1'h0)] wire215;
  wire signed [(5'h12):(1'h0)] wire79;
  wire [(4'hb):(1'h0)] wire78;
  wire signed [(5'h11):(1'h0)] wire77;
  wire signed [(3'h4):(1'h0)] wire76;
  reg signed [(4'he):(1'h0)] reg75 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg74 = (1'h0);
  reg signed [(4'he):(1'h0)] reg73 = (1'h0);
  reg [(5'h15):(1'h0)] reg72 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg71 = (1'h0);
  reg [(3'h6):(1'h0)] reg70 = (1'h0);
  reg [(5'h11):(1'h0)] reg69 = (1'h0);
  reg [(3'h7):(1'h0)] reg68 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg67 = (1'h0);
  reg [(5'h14):(1'h0)] reg66 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg65 = (1'h0);
  reg [(5'h10):(1'h0)] reg64 = (1'h0);
  reg [(5'h15):(1'h0)] reg63 = (1'h0);
  reg [(4'hf):(1'h0)] reg62 = (1'h0);
  reg [(3'h6):(1'h0)] reg61 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg60 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire59;
  wire signed [(4'he):(1'h0)] wire58;
  wire [(5'h11):(1'h0)] wire57;
  reg [(5'h15):(1'h0)] reg56 = (1'h0);
  reg [(3'h6):(1'h0)] reg55 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg54 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg53 = (1'h0);
  reg [(4'h9):(1'h0)] reg52 = (1'h0);
  reg [(4'h9):(1'h0)] reg51 = (1'h0);
  reg [(5'h10):(1'h0)] reg50 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg49 = (1'h0);
  wire [(4'hb):(1'h0)] wire48;
  reg [(4'he):(1'h0)] reg47 = (1'h0);
  wire [(5'h14):(1'h0)] wire45;
  wire signed [(5'h15):(1'h0)] wire217;
  wire [(2'h2):(1'h0)] wire218;
  assign y = {reg226,
                 reg225,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 wire215,
                 wire79,
                 wire78,
                 wire77,
                 wire76,
                 reg75,
                 reg74,
                 reg73,
                 reg72,
                 reg71,
                 reg70,
                 reg69,
                 reg68,
                 reg67,
                 reg66,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 wire59,
                 wire58,
                 wire57,
                 reg56,
                 reg55,
                 reg54,
                 reg53,
                 reg52,
                 reg51,
                 reg50,
                 reg49,
                 wire48,
                 reg47,
                 wire45,
                 wire217,
                 wire218,
                 (1'h0)};
  module4 modinst46 (.wire7(wire3), .wire5(wire2), .wire8(wire0), .wire6(wire1), .y(wire45), .clk(clk));
  always
    @(posedge clk) begin
      reg47 <= wire3[(4'hc):(4'ha)];
    end
  assign wire48 = $unsigned($signed({$unsigned($signed((8'ha8))),
                      ((wire45 <<< wire1) < $signed((8'haf)))}));
  always
    @(posedge clk) begin
      if (wire1)
        begin
          reg49 <= ($unsigned((wire3 ?
              wire0[(4'h8):(3'h5)] : ((wire0 ?
                  wire48 : wire0) ^ wire2[(3'h6):(3'h5)]))) >= wire3);
          reg50 <= {(~^(wire1 ? $unsigned($unsigned(wire48)) : wire48)),
              (wire1 ?
                  ({(-wire0),
                      (8'hbd)} + reg47[(4'ha):(1'h0)]) : ((wire1[(1'h0):(1'h0)] ?
                          wire2 : wire1[(2'h2):(1'h1)]) ?
                      wire0 : wire48))};
          reg51 <= $unsigned({{($signed(reg49) ^ wire1[(4'hc):(4'hb)]),
                  reg49[(1'h0):(1'h0)]},
              (((reg47 - wire3) ?
                  (wire45 ?
                      wire2 : wire2) : (|wire1)) >> wire0[(4'ha):(4'h9)])});
        end
      else
        begin
          reg49 <= $unsigned((wire48 ^ (~|($signed((8'hb6)) && (~wire1)))));
          reg50 <= $unsigned((~&{wire2}));
          if (((($unsigned(wire45[(4'h8):(3'h5)]) ? wire0 : {(7'h41)}) ?
                  (($signed(reg51) >>> (wire45 != reg51)) ?
                      (((8'ha4) ? wire48 : wire45) ?
                          reg47 : reg51[(4'h9):(1'h1)]) : $unsigned((8'hbf))) : ($unsigned($unsigned(wire45)) == $signed(reg49))) ?
              (^~(8'hac)) : reg50))
            begin
              reg51 <= wire2;
              reg52 <= $signed((reg47[(4'hc):(4'h9)] >> wire2));
              reg53 <= (8'hab);
              reg54 <= (({wire48} ?
                  $unsigned($signed((~wire3))) : {(7'h44)}) >>> ((&(wire45 | (wire1 ^ reg51))) & reg51[(2'h3):(1'h1)]));
              reg55 <= ((~|((reg53 & wire45[(5'h14):(5'h10)]) ?
                  $signed($unsigned(reg51)) : wire48)) >= $unsigned((8'hb8)));
            end
          else
            begin
              reg51 <= (((reg55 ~^ {$unsigned((8'ha8)), $unsigned(reg52)}) ?
                  reg50[(3'h6):(1'h1)] : $signed((+wire0))) ^~ (8'ha1));
              reg52 <= reg54;
              reg53 <= $signed(wire3);
              reg54 <= $signed(({$signed((^wire3))} <= wire45));
            end
          reg56 <= wire45[(3'h7):(1'h1)];
        end
    end
  assign wire57 = $unsigned($unsigned((!$signed((+(7'h42))))));
  assign wire58 = (!wire3[(2'h2):(1'h1)]);
  assign wire59 = reg47;
  always
    @(posedge clk) begin
      reg60 <= wire0[(3'h6):(2'h3)];
      if ($signed(wire59[(4'hd):(3'h4)]))
        begin
          if (($unsigned(reg50) >> wire48))
            begin
              reg61 <= wire57;
              reg62 <= reg55[(2'h3):(1'h0)];
              reg63 <= {$signed(wire57[(1'h0):(1'h0)])};
            end
          else
            begin
              reg61 <= wire3;
              reg62 <= $signed($signed(reg49));
            end
          reg64 <= wire0[(2'h2):(1'h0)];
        end
      else
        begin
          reg61 <= (($unsigned({$signed(reg55), $signed(wire59)}) ?
                  reg64 : {reg56[(4'ha):(3'h4)], reg56}) ?
              ($signed(({reg54,
                  wire59} ^~ wire48[(4'h8):(2'h3)])) ^ (-((~&reg64) ?
                  (wire2 != reg56) : {wire45, wire3}))) : ($unsigned(wire58) ?
                  {$unsigned(wire59)} : $signed(((reg55 >= reg47) ^ (wire48 - reg62)))));
          if (reg54)
            begin
              reg62 <= $unsigned($unsigned((+((^~(8'hb6)) ?
                  wire45 : $unsigned(reg49)))));
            end
          else
            begin
              reg62 <= reg56;
              reg63 <= (reg60[(2'h3):(1'h0)] > (!(wire58[(4'h9):(4'h8)] << (((8'hb2) & wire45) & (wire3 == reg50)))));
              reg64 <= ({(((reg52 >>> reg49) ? (wire3 - reg64) : (+(8'hb7))) ?
                          reg64[(3'h4):(3'h4)] : $unsigned((reg51 ?
                              reg47 : reg54)))} ?
                  {($unsigned(wire48[(3'h7):(3'h7)]) ?
                          {wire3[(3'h4):(1'h0)],
                              $unsigned(reg54)} : reg61)} : wire2);
              reg65 <= (reg52[(3'h6):(3'h4)] ?
                  (-(reg60[(3'h5):(2'h3)] ?
                      reg49[(4'hb):(4'ha)] : $signed(wire3))) : {(((reg62 | reg50) ?
                          $unsigned(reg60) : $unsigned((8'hbf))) * ((~wire48) ?
                          reg60 : (wire59 ? wire0 : wire2))),
                      $unsigned($unsigned((+reg55)))});
            end
          reg66 <= ({(($signed(reg64) ?
                          $unsigned(wire0) : wire1[(4'ha):(3'h6)]) ?
                      (~$unsigned((7'h41))) : (^(+wire58)))} ?
              reg63[(3'h7):(3'h4)] : (($signed($signed(reg61)) <= $signed($signed((8'had)))) >> wire59[(4'ha):(2'h3)]));
          reg67 <= ($signed($unsigned({(reg65 ? wire59 : reg49)})) ?
              wire59[(4'hd):(4'hb)] : ((~^($unsigned(wire3) ? reg53 : wire3)) ?
                  $unsigned(($unsigned(wire48) < $unsigned(wire3))) : $unsigned(($unsigned(reg49) ?
                      reg49[(2'h2):(1'h0)] : (reg61 - (8'hb6))))));
          reg68 <= ((wire2[(2'h2):(2'h2)] ?
                  ($unsigned((^reg61)) ?
                      (8'hb5) : $signed(reg61[(1'h1):(1'h0)])) : ($signed($unsigned(wire57)) <= reg53[(4'h8):(3'h7)])) ?
              ($unsigned(wire59) != wire1) : $unsigned(reg49));
        end
      if ((^~(reg54[(2'h3):(2'h3)] ?
          (reg47 > reg56) : $unsigned($signed($unsigned(reg67))))))
        begin
          reg69 <= reg53[(3'h5):(1'h0)];
          reg70 <= reg52;
          reg71 <= $unsigned({$signed(((wire48 * reg63) ? reg53 : {reg47})),
              (reg62[(3'h4):(2'h3)] ? {wire45, wire57} : $signed((~|wire48)))});
          reg72 <= wire57;
          reg73 <= reg64[(5'h10):(1'h1)];
        end
      else
        begin
          reg69 <= ($signed((wire0 ?
                  ($unsigned(reg73) ? {reg70} : wire48) : {reg53[(3'h4):(2'h2)],
                      (&wire0)})) ?
              ((~^(-(|reg49))) >> (($unsigned(wire58) ?
                  $unsigned(reg70) : {reg61,
                      wire48}) ^~ $signed((reg54 <= reg71)))) : reg52);
          if (((reg50[(4'hc):(1'h1)] == reg53) < reg70))
            begin
              reg70 <= {wire2[(3'h5):(1'h0)]};
              reg71 <= wire2[(4'h8):(3'h4)];
              reg72 <= {reg51};
            end
          else
            begin
              reg70 <= {wire3};
            end
          reg73 <= $signed(reg70[(1'h1):(1'h0)]);
          reg74 <= reg52;
          reg75 <= reg68[(2'h2):(1'h1)];
        end
    end
  assign wire76 = $unsigned((~^reg66));
  assign wire77 = (reg73 << $unsigned((~({wire76} || (reg64 ?
                      reg61 : wire48)))));
  assign wire78 = (8'haa);
  assign wire79 = reg64;
  module80 modinst216 (wire215, clk, reg69, reg72, wire2, reg50, wire0);
  assign wire217 = {reg64};
  module13 modinst219 (wire218, clk, wire217, reg52, wire0, wire2, wire57);
  always
    @(posedge clk) begin
      reg220 <= (7'h40);
      reg221 <= $signed(($unsigned((reg47[(3'h5):(2'h3)] | (^(8'hb3)))) ?
          ({reg65[(2'h3):(2'h3)], reg56[(5'h12):(4'h9)]} + ((wire45 ?
                  reg49 : wire218) ?
              (reg55 ?
                  (8'h9f) : reg50) : $signed(reg53))) : ($unsigned((wire78 ?
                  wire217 : reg68)) ?
              $unsigned(wire3[(4'h9):(2'h3)]) : (~&reg50))));
      if (((($signed($unsigned(reg70)) - $unsigned((reg61 <<< reg47))) > (8'hab)) ?
          ($unsigned($unsigned($signed((8'hbb)))) ?
              (-wire218) : (8'ha7)) : $signed(wire1)))
        begin
          if ((&$unsigned((reg221 | {{(8'hba)}}))))
            begin
              reg222 <= wire218;
            end
          else
            begin
              reg222 <= $signed((|$signed(wire48)));
              reg223 <= {$unsigned(($unsigned($signed(reg75)) ~^ wire78)),
                  reg71};
              reg224 <= (8'hbb);
            end
          reg225 <= $unsigned(wire58);
          reg226 <= (~|reg74[(4'hf):(4'hf)]);
        end
      else
        begin
          reg222 <= reg66;
          reg223 <= ($unsigned($signed(reg63[(3'h7):(2'h2)])) ?
              (^wire59) : reg223[(1'h1):(1'h0)]);
        end
    end
endmodule

module module80
#( parameter param214 = (~|(~|((((8'hac) << (8'ha5)) > ((8'hb5) > (8'haa))) ? (((8'hbc) > (8'h9c)) ? ((8'hbc) > (8'ha4)) : (~|(8'ha0))) : ({(7'h41), (7'h40)} ? ((8'h9e) ? (8'hb6) : (8'hbe)) : (~(8'ha8)))))) )
(y, clk, wire81, wire82, wire83, wire84, wire85);
  output wire [(32'ha2):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire81;
  input wire [(3'h7):(1'h0)] wire82;
  input wire signed [(4'ha):(1'h0)] wire83;
  input wire [(3'h6):(1'h0)] wire84;
  input wire signed [(5'h13):(1'h0)] wire85;
  wire signed [(2'h3):(1'h0)] wire213;
  wire [(2'h2):(1'h0)] wire212;
  wire signed [(5'h15):(1'h0)] wire210;
  wire signed [(4'hf):(1'h0)] wire176;
  wire [(3'h4):(1'h0)] wire86;
  wire [(3'h5):(1'h0)] wire87;
  wire [(4'hb):(1'h0)] wire88;
  reg [(5'h11):(1'h0)] reg89 = (1'h0);
  wire [(5'h12):(1'h0)] wire90;
  wire [(4'hb):(1'h0)] wire91;
  wire signed [(4'h8):(1'h0)] wire92;
  wire [(3'h5):(1'h0)] wire93;
  wire [(5'h14):(1'h0)] wire94;
  wire signed [(5'h15):(1'h0)] wire174;
  assign y = {wire213,
                 wire212,
                 wire210,
                 wire176,
                 wire86,
                 wire87,
                 wire88,
                 reg89,
                 wire90,
                 wire91,
                 wire92,
                 wire93,
                 wire94,
                 wire174,
                 (1'h0)};
  assign wire86 = (^~(wire85[(2'h2):(2'h2)] ?
                      $unsigned(($unsigned(wire84) | (wire81 != wire83))) : (^{wire83})));
  assign wire87 = wire83;
  assign wire88 = (8'hac);
  always
    @(posedge clk) begin
      reg89 <= (|(wire81 != (($signed(wire83) ?
          (wire87 ? wire88 : (8'ha9)) : (wire87 ?
              wire83 : (8'ha5))) << (~(~|wire87)))));
    end
  assign wire90 = $unsigned((&($signed($unsigned(reg89)) >>> ((^~wire83) < $unsigned((8'ha3))))));
  assign wire91 = wire82[(3'h7):(3'h5)];
  assign wire92 = (($signed(($unsigned(wire86) ?
                      reg89[(2'h2):(1'h0)] : $unsigned(wire81))) && wire91[(4'h8):(4'h8)]) < {wire83,
                      (wire86 | ($signed(wire91) ?
                          $unsigned(wire88) : (wire82 ? wire85 : wire87)))});
  assign wire93 = wire92[(3'h6):(3'h4)];
  assign wire94 = ((-(^{(^~wire91)})) << wire92[(3'h4):(2'h3)]);
  module95 modinst175 (.y(wire174), .wire97(wire94), .clk(clk), .wire98(wire88), .wire100(wire83), .wire96(reg89), .wire99(wire86));
  assign wire176 = (-(^~$unsigned(wire85[(2'h2):(2'h2)])));
  module177 modinst211 (.y(wire210), .wire180(wire84), .wire181(wire85), .wire179(wire82), .wire178(wire81), .clk(clk));
  assign wire212 = (wire85 - ((!wire82[(3'h5):(3'h4)]) ~^ ($signed((wire81 || wire210)) ?
                       $unsigned($unsigned(wire87)) : wire86)));
  assign wire213 = wire88;
endmodule

module module4  (y, clk, wire8, wire7, wire6, wire5);
  output wire [(32'h8b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h7):(1'h0)] wire8;
  input wire [(5'h11):(1'h0)] wire7;
  input wire [(4'hc):(1'h0)] wire6;
  input wire [(4'hb):(1'h0)] wire5;
  wire signed [(4'hd):(1'h0)] wire44;
  wire signed [(2'h2):(1'h0)] wire43;
  wire signed [(5'h11):(1'h0)] wire42;
  wire signed [(5'h11):(1'h0)] wire24;
  wire signed [(5'h12):(1'h0)] wire12;
  wire signed [(5'h14):(1'h0)] wire11;
  wire signed [(5'h13):(1'h0)] wire10;
  wire [(5'h14):(1'h0)] wire9;
  wire [(4'hc):(1'h0)] wire40;
  assign y = {wire44,
                 wire43,
                 wire42,
                 wire24,
                 wire12,
                 wire11,
                 wire10,
                 wire9,
                 wire40,
                 (1'h0)};
  assign wire9 = $unsigned((wire8[(2'h2):(1'h1)] + $unsigned($signed($unsigned(wire7)))));
  assign wire10 = (&(~|(wire5[(1'h0):(1'h0)] ?
                      wire6[(4'hc):(2'h3)] : (((8'hb5) >>> (8'haa)) | (wire8 ?
                          wire7 : wire6)))));
  assign wire11 = ($signed(wire6) != (!($unsigned((wire8 >= wire8)) ^ wire9)));
  assign wire12 = ($unsigned({{wire5[(4'h9):(3'h7)]}, wire6}) ?
                      (8'hae) : (~&wire10[(4'hd):(4'hd)]));
  module13 modinst25 (.wire16(wire11), .wire15(wire9), .wire18(wire10), .clk(clk), .wire14(wire7), .y(wire24), .wire17(wire12));
  module26 modinst41 (wire40, clk, wire10, wire24, wire5, wire11, wire12);
  assign wire42 = (+$unsigned($unsigned(wire40)));
  assign wire43 = ((|({$signed(wire11)} | wire10[(4'hf):(3'h5)])) ?
                      (wire42 ?
                          ($unsigned({wire9,
                              wire11}) | $signed($signed(wire7))) : wire6[(3'h5):(1'h0)]) : ((+$unsigned(wire5)) >> {((wire5 ?
                              (8'hac) : wire11) & (-wire24)),
                          (+$signed((7'h43)))}));
  assign wire44 = $signed((~&(~^{$signed(wire43)})));
endmodule

module module26
#( parameter param38 = ((((((7'h44) + (8'hb9)) >> ((8'ha3) ~^ (8'h9c))) ? (((8'hb6) ? (8'hbc) : (7'h43)) ~^ ((7'h43) >= (8'hbb))) : {(&(8'hb7))}) & ((8'hb1) ? ((~&(8'ha1)) ? {(8'ha8), (8'ha0)} : (7'h41)) : {((7'h44) ? (8'h9d) : (7'h42))})) ? (|((&(^~(8'had))) <= (~&(~&(8'ha8))))) : ((+{((8'haa) ? (8'hbb) : (8'h9d))}) ? ((((8'ha1) ? (8'ha6) : (8'had)) ? (~&(7'h42)) : (-(8'ha5))) == {(~|(8'ha8))}) : (({(8'ha7), (8'haa)} << (~|(8'ha9))) <<< ({(8'hb9), (8'hbd)} - {(7'h41)}))))
, parameter param39 = (({((param38 ? param38 : param38) ? (param38 >>> param38) : (param38 ? param38 : param38)), (^~{param38, param38})} && param38) ? param38 : ({(param38 < (param38 * param38))} ? (~{{param38, (8'hab)}, param38}) : {(&(param38 ? (7'h43) : param38)), (~(param38 ? param38 : param38))})) )
(y, clk, wire31, wire30, wire29, wire28, wire27);
  output wire [(32'h4b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire31;
  input wire [(3'h4):(1'h0)] wire30;
  input wire [(3'h7):(1'h0)] wire29;
  input wire [(5'h14):(1'h0)] wire28;
  input wire [(5'h12):(1'h0)] wire27;
  wire [(4'hc):(1'h0)] wire37;
  wire [(4'h9):(1'h0)] wire36;
  wire signed [(5'h15):(1'h0)] wire35;
  wire [(4'he):(1'h0)] wire34;
  wire [(2'h3):(1'h0)] wire33;
  wire [(4'hf):(1'h0)] wire32;
  assign y = {wire37, wire36, wire35, wire34, wire33, wire32, (1'h0)};
  assign wire32 = (($unsigned($signed($signed(wire28))) * ((!{wire28}) && (&(wire31 | wire31)))) ?
                      (({{wire27}} ^ ($unsigned(wire28) <= {wire31, wire27})) ?
                          ($signed(wire31[(3'h6):(3'h6)]) ?
                              ((wire29 ?
                                  wire28 : wire27) << wire27) : (~|(wire31 << wire28))) : ($signed($signed(wire28)) ?
                              wire30 : ($unsigned(wire29) ?
                                  wire28 : (wire27 ^~ wire31)))) : $signed({{$signed(wire28)}}));
  assign wire33 = (wire28[(3'h7):(3'h7)] == (($signed((|(7'h44))) ~^ $signed((wire32 > wire32))) > $unsigned($signed($unsigned(wire29)))));
  assign wire34 = wire32[(4'hc):(1'h0)];
  assign wire35 = $signed((^~$signed(wire33)));
  assign wire36 = ((~&$signed(wire31)) * ((({wire29} && (wire29 & wire28)) & $unsigned(wire29)) << (^((wire31 ^ wire33) ?
                      {wire29, wire33} : ((8'ha9) ? wire34 : wire29)))));
  assign wire37 = wire34[(3'h6):(3'h5)];
endmodule

module module13
#( parameter param23 = {(((~((8'h9f) ? (8'ha8) : (8'hab))) * (7'h42)) || {(((8'hb1) < (8'haf)) <= ((8'h9d) ? (8'had) : (8'hba))), (((8'ha5) ? (8'hbf) : (7'h42)) * ((8'h9c) > (7'h44)))}), {(&(((8'ha1) ? (8'ha8) : (8'hb4)) ? ((8'hb6) ? (8'hbc) : (8'hb1)) : {(8'hb5)}))}} )
(y, clk, wire18, wire17, wire16, wire15, wire14);
  output wire [(32'h43):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h13):(1'h0)] wire18;
  input wire signed [(4'h9):(1'h0)] wire17;
  input wire [(4'hf):(1'h0)] wire16;
  input wire [(5'h14):(1'h0)] wire15;
  input wire [(5'h11):(1'h0)] wire14;
  wire [(4'hc):(1'h0)] wire22;
  wire signed [(5'h14):(1'h0)] wire21;
  wire signed [(5'h14):(1'h0)] wire20;
  reg [(4'he):(1'h0)] reg19 = (1'h0);
  assign y = {wire22, wire21, wire20, reg19, (1'h0)};
  always
    @(posedge clk) begin
      reg19 <= $signed(wire17);
    end
  assign wire20 = ((wire15[(5'h12):(5'h12)] >>> $signed(((wire18 << wire14) <= $signed(wire17)))) * $signed(((~&$unsigned(wire18)) ?
                      ($unsigned(reg19) ?
                          (wire17 < wire15) : (~|(8'hb7))) : {(wire14 ?
                              reg19 : wire16)})));
  assign wire21 = (+((~|$signed(wire17[(3'h5):(3'h5)])) ^ (+({wire17,
                      wire14} < wire18))));
  assign wire22 = (-$unsigned((wire17 * {$unsigned(reg19), {wire17}})));
endmodule

module module177  (y, clk, wire181, wire180, wire179, wire178);
  output wire [(32'h12f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire181;
  input wire signed [(3'h5):(1'h0)] wire180;
  input wire [(2'h3):(1'h0)] wire179;
  input wire [(4'ha):(1'h0)] wire178;
  wire [(5'h11):(1'h0)] wire209;
  wire signed [(5'h14):(1'h0)] wire208;
  wire signed [(4'hc):(1'h0)] wire207;
  wire [(5'h13):(1'h0)] wire206;
  wire [(3'h7):(1'h0)] wire205;
  wire signed [(3'h4):(1'h0)] wire204;
  wire [(5'h13):(1'h0)] wire203;
  reg signed [(3'h7):(1'h0)] reg202 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg201 = (1'h0);
  reg [(3'h4):(1'h0)] reg200 = (1'h0);
  reg [(5'h11):(1'h0)] reg199 = (1'h0);
  reg [(4'hb):(1'h0)] reg198 = (1'h0);
  reg [(4'hf):(1'h0)] reg197 = (1'h0);
  reg [(5'h15):(1'h0)] reg196 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire195;
  wire signed [(3'h6):(1'h0)] wire194;
  wire signed [(5'h13):(1'h0)] wire193;
  wire [(4'hb):(1'h0)] wire192;
  wire signed [(4'hf):(1'h0)] wire191;
  wire signed [(4'hb):(1'h0)] wire190;
  wire [(2'h3):(1'h0)] wire189;
  wire [(4'hc):(1'h0)] wire188;
  wire signed [(5'h10):(1'h0)] wire187;
  wire signed [(2'h3):(1'h0)] wire186;
  wire signed [(3'h4):(1'h0)] wire185;
  wire signed [(2'h3):(1'h0)] wire184;
  wire [(4'ha):(1'h0)] wire183;
  reg signed [(4'h9):(1'h0)] reg182 = (1'h0);
  assign y = {wire209,
                 wire208,
                 wire207,
                 wire206,
                 wire205,
                 wire204,
                 wire203,
                 reg202,
                 reg201,
                 reg200,
                 reg199,
                 reg198,
                 reg197,
                 reg196,
                 wire195,
                 wire194,
                 wire193,
                 wire192,
                 wire191,
                 wire190,
                 wire189,
                 wire188,
                 wire187,
                 wire186,
                 wire185,
                 wire184,
                 wire183,
                 reg182,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg182 <= wire179[(1'h1):(1'h1)];
    end
  assign wire183 = $signed($unsigned({($unsigned(wire180) << wire181),
                       $unsigned($unsigned((8'ha6)))}));
  assign wire184 = (+wire181[(5'h10):(4'hf)]);
  assign wire185 = {$unsigned(wire178), $signed(wire178[(4'ha):(3'h6)])};
  assign wire186 = $unsigned({wire179[(2'h2):(1'h0)],
                       (^wire180[(3'h5):(3'h4)])});
  assign wire187 = $signed((~^(wire180 ?
                       $unsigned(wire183) : ({wire178,
                           reg182} << wire184[(1'h0):(1'h0)]))));
  assign wire188 = $signed(((($signed(wire185) ?
                       {(8'ha1), wire181} : (8'h9d)) <= $signed((wire185 ?
                       wire183 : wire179))) ~^ $signed((|(wire181 ?
                       wire186 : wire185)))));
  assign wire189 = $unsigned(($signed(wire185) ?
                       $unsigned((~^$unsigned(wire188))) : $signed(wire178)));
  assign wire190 = (7'h44);
  assign wire191 = {$unsigned($signed((wire179[(2'h2):(2'h2)] | {wire181,
                           wire179})))};
  assign wire192 = $unsigned((~|$unsigned(wire189[(2'h3):(1'h1)])));
  assign wire193 = ((($unsigned($unsigned(wire187)) + $signed(wire191[(4'hd):(1'h0)])) ?
                           $unsigned({wire178[(2'h2):(1'h0)]}) : $signed((^~$unsigned(wire192)))) ?
                       {$signed((~&(wire183 ? wire185 : wire180))),
                           wire179[(1'h1):(1'h0)]} : ({((wire186 || wire185) <<< (wire186 ?
                                   wire191 : (8'hab))),
                               $signed($unsigned(wire187))} ?
                           (~|wire178[(4'h9):(3'h5)]) : wire191));
  assign wire194 = (^wire188[(2'h2):(2'h2)]);
  assign wire195 = {(!(reg182 ? wire188 : wire194)),
                       ($signed(({wire187, wire190} ?
                           $unsigned(reg182) : $signed(wire183))) & $unsigned($signed((wire192 ?
                           wire189 : wire184))))};
  always
    @(posedge clk) begin
      reg196 <= $signed(wire185[(2'h2):(1'h1)]);
      reg197 <= $signed(reg182[(3'h7):(1'h0)]);
      if ($unsigned($unsigned(wire183[(1'h0):(1'h0)])))
        begin
          reg198 <= (!$unsigned($unsigned(wire186[(2'h2):(1'h1)])));
          reg199 <= $unsigned({$signed((~|(wire178 ? wire178 : wire188)))});
          if (({{wire183,
                  {$unsigned(reg197)}}} == $unsigned($signed($signed((wire192 ?
              wire193 : (8'ha0)))))))
            begin
              reg200 <= ((~|reg197) ?
                  $unsigned((~&$unsigned(wire178[(4'ha):(4'h9)]))) : reg198);
              reg201 <= wire191;
            end
          else
            begin
              reg200 <= wire178;
              reg201 <= (~(wire186 ?
                  $unsigned(((reg199 | wire189) ^ ((8'hb5) >> wire178))) : (8'h9d)));
            end
        end
      else
        begin
          reg198 <= (8'hac);
          reg199 <= (($signed(reg197) && $unsigned((~^(~(8'ha2))))) ~^ $unsigned(($signed((wire183 ~^ (8'ha0))) ?
              ($unsigned(reg198) ?
                  (&(8'ha4)) : (wire192 ?
                      (7'h42) : wire189)) : (wire184[(1'h1):(1'h0)] & $unsigned(wire190)))));
          reg200 <= ($signed(wire180) | (^wire195));
        end
      reg202 <= ((~|reg196[(4'h8):(3'h6)]) ~^ (wire187[(3'h5):(1'h1)] != (($unsigned(wire188) ?
              (+wire190) : wire189) ?
          reg196[(4'hc):(3'h7)] : {$unsigned(wire193), (wire190 || (8'hbe))})));
    end
  assign wire203 = ((8'hb3) ?
                       {{({wire184} ?
                                   wire180[(3'h4):(2'h2)] : $signed(reg200))},
                           reg196[(4'ha):(4'h9)]} : (+wire193));
  assign wire204 = (-reg201);
  assign wire205 = wire181[(4'ha):(2'h3)];
  assign wire206 = {$signed(wire186), wire193[(4'h9):(1'h0)]};
  assign wire207 = reg197[(2'h3):(1'h1)];
  assign wire208 = $signed($signed($signed($signed({wire195, wire180}))));
  assign wire209 = ((~&({((8'hb0) ? wire194 : reg198),
                           (wire208 > wire192)} >> (^$unsigned(wire180)))) ?
                       (^~$signed(($unsigned(wire206) - (wire206 ?
                           (8'haf) : wire207)))) : $unsigned(((!(+reg196)) ?
                           ($signed(wire185) == (^wire205)) : (~&wire206))));
endmodule

module module95
#( parameter param173 = ((8'h9f) ? ((({(8'ha2), (8'ha5)} ? {(8'hab), (8'hb9)} : (+(8'hb4))) | ((~&(8'had)) ? ((8'hb7) ^ (7'h44)) : (&(8'ha0)))) ? (-{(-(8'ha3))}) : (8'hab)) : (^~(&((~(8'hb6)) <<< ((8'hab) > (8'hb8)))))) )
(y, clk, wire100, wire99, wire98, wire97, wire96);
  output wire [(32'h33c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire100;
  input wire [(3'h4):(1'h0)] wire99;
  input wire signed [(2'h2):(1'h0)] wire98;
  input wire [(2'h2):(1'h0)] wire97;
  input wire [(4'hf):(1'h0)] wire96;
  reg signed [(4'h8):(1'h0)] reg172 = (1'h0);
  reg [(4'hd):(1'h0)] reg171 = (1'h0);
  reg [(5'h12):(1'h0)] reg170 = (1'h0);
  reg [(4'hd):(1'h0)] reg169 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg168 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg167 = (1'h0);
  reg [(5'h15):(1'h0)] reg166 = (1'h0);
  reg [(2'h3):(1'h0)] reg165 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg164 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg163 = (1'h0);
  reg [(4'hc):(1'h0)] reg162 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg161 = (1'h0);
  reg [(4'he):(1'h0)] reg160 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg159 = (1'h0);
  reg [(4'h9):(1'h0)] reg158 = (1'h0);
  reg [(3'h6):(1'h0)] reg157 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg156 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg155 = (1'h0);
  reg [(4'hf):(1'h0)] reg154 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg153 = (1'h0);
  reg [(5'h14):(1'h0)] reg152 = (1'h0);
  reg [(5'h10):(1'h0)] reg151 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg150 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg149 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg148 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg147 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg146 = (1'h0);
  reg [(4'h9):(1'h0)] reg145 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg144 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire143;
  reg [(4'h8):(1'h0)] reg142 = (1'h0);
  reg [(4'h8):(1'h0)] reg141 = (1'h0);
  reg [(5'h15):(1'h0)] reg140 = (1'h0);
  reg [(4'hc):(1'h0)] reg139 = (1'h0);
  reg [(5'h15):(1'h0)] reg138 = (1'h0);
  wire [(3'h7):(1'h0)] wire137;
  wire [(3'h4):(1'h0)] wire136;
  reg [(4'hd):(1'h0)] reg135 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg134 = (1'h0);
  reg [(2'h3):(1'h0)] reg133 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg132 = (1'h0);
  reg [(4'hb):(1'h0)] reg131 = (1'h0);
  reg [(5'h11):(1'h0)] reg130 = (1'h0);
  reg [(3'h6):(1'h0)] reg129 = (1'h0);
  reg [(3'h6):(1'h0)] reg128 = (1'h0);
  reg [(3'h6):(1'h0)] reg127 = (1'h0);
  wire [(4'h9):(1'h0)] wire126;
  wire [(4'he):(1'h0)] wire125;
  reg [(5'h15):(1'h0)] reg124 = (1'h0);
  reg [(4'hd):(1'h0)] reg123 = (1'h0);
  reg [(4'ha):(1'h0)] reg122 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg121 = (1'h0);
  reg [(4'hd):(1'h0)] reg120 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg119 = (1'h0);
  reg [(2'h3):(1'h0)] reg118 = (1'h0);
  reg [(4'h9):(1'h0)] reg117 = (1'h0);
  reg [(4'hb):(1'h0)] reg116 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg115 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg114 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg113 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg112 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg111 = (1'h0);
  reg [(4'he):(1'h0)] reg110 = (1'h0);
  reg [(4'hf):(1'h0)] reg109 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg108 = (1'h0);
  reg [(5'h15):(1'h0)] reg107 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg106 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg105 = (1'h0);
  reg [(4'h9):(1'h0)] reg104 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg103 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg102 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire101;
  assign y = {reg172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 reg149,
                 reg148,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 wire143,
                 reg142,
                 reg141,
                 reg140,
                 reg139,
                 reg138,
                 wire137,
                 wire136,
                 reg135,
                 reg134,
                 reg133,
                 reg132,
                 reg131,
                 reg130,
                 reg129,
                 reg128,
                 reg127,
                 wire126,
                 wire125,
                 reg124,
                 reg123,
                 reg122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 reg117,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 reg112,
                 reg111,
                 reg110,
                 reg109,
                 reg108,
                 reg107,
                 reg106,
                 reg105,
                 reg104,
                 reg103,
                 reg102,
                 wire101,
                 (1'h0)};
  assign wire101 = {$signed((~|wire96[(3'h4):(1'h0)])), wire100};
  always
    @(posedge clk) begin
      if (wire99)
        begin
          reg102 <= (wire100[(4'h9):(4'h9)] ?
              $unsigned(($signed(wire97[(1'h0):(1'h0)]) ?
                  ((wire100 != wire96) ?
                      {wire101,
                          (8'ha6)} : (|wire97)) : $unsigned($signed(wire99)))) : (&(wire100[(1'h0):(1'h0)] ^~ (&(wire101 ?
                  (8'had) : wire97)))));
        end
      else
        begin
          reg102 <= $signed(wire101);
          reg103 <= wire101[(1'h1):(1'h0)];
          reg104 <= $signed((reg102[(1'h0):(1'h0)] ?
              ((|((8'haf) << wire96)) ?
                  $signed((wire98 ? wire97 : reg103)) : $unsigned((reg102 ?
                      wire98 : wire100))) : wire97));
          reg105 <= reg104[(3'h7):(1'h0)];
          reg106 <= $unsigned(wire100);
        end
      reg107 <= (8'ha2);
      if (($unsigned(wire98) && wire97[(1'h0):(1'h0)]))
        begin
          reg108 <= ($unsigned(reg107) && (+(reg106 - $signed((wire97 || wire101)))));
          reg109 <= (~wire97);
          reg110 <= (~^$unsigned((^$signed((reg107 ~^ wire98)))));
          reg111 <= reg104;
        end
      else
        begin
          if ($unsigned((wire97[(2'h2):(1'h1)] ^~ (reg110[(3'h6):(3'h6)] <<< $signed(wire98)))))
            begin
              reg108 <= {({$unsigned($signed((7'h42))),
                      wire99} && $signed(wire101)),
                  $unsigned(wire98)};
            end
          else
            begin
              reg108 <= $unsigned((reg106[(4'h8):(2'h2)] ?
                  wire99[(1'h1):(1'h1)] : (~(reg108 ?
                      $unsigned(reg111) : (reg107 ? reg109 : reg104)))));
              reg109 <= wire97;
              reg110 <= wire100;
              reg111 <= (8'hb5);
            end
          if ((({reg105[(3'h7):(3'h7)], reg109[(3'h6):(1'h1)]} || (~&(reg104 ?
              reg105[(3'h7):(3'h5)] : (+(8'ha2))))) & {{(8'ha3), reg110}}))
            begin
              reg112 <= $signed((8'haf));
              reg113 <= wire100;
              reg114 <= reg103;
              reg115 <= reg110;
              reg116 <= wire97[(1'h0):(1'h0)];
            end
          else
            begin
              reg112 <= $unsigned((~|(!($unsigned(wire97) || reg105[(3'h7):(1'h0)]))));
            end
          if ({(($signed(reg111) <= (~|(reg110 >>> reg114))) == wire96[(3'h4):(2'h2)]),
              reg104})
            begin
              reg117 <= $unsigned(($unsigned((~&(^(8'hb5)))) >> (reg103 ?
                  ({reg106,
                      reg114} * wire100[(2'h2):(2'h2)]) : $signed(wire96[(1'h1):(1'h1)]))));
              reg118 <= ((8'hb3) ?
                  reg109 : ({wire101, $signed((&reg105))} ^ reg103));
            end
          else
            begin
              reg117 <= ((^~($unsigned(reg116) - ((+reg116) - reg104[(2'h2):(2'h2)]))) ^~ ((($signed((8'hb0)) ?
                          (~wire98) : {wire96}) ?
                      $unsigned(wire96[(4'h9):(3'h6)]) : $signed(reg114)) ?
                  $unsigned({(reg115 + wire97),
                      (reg112 ? reg105 : wire96)}) : ((wire97 ?
                          wire100[(3'h7):(1'h0)] : $signed(reg118)) ?
                      $signed((+reg108)) : (~|(reg109 ? reg102 : wire101)))));
            end
          if ((((($unsigned((8'h9d)) ^~ ((8'hbf) ?
                      wire96 : wire96)) != wire96) ?
                  (reg117 != (|(!reg110))) : reg117[(4'h8):(3'h5)]) ?
              (^~(8'hae)) : ((reg110 == (reg117 < {reg118})) + $signed($unsigned($signed(reg117))))))
            begin
              reg119 <= $signed(reg115);
              reg120 <= {(reg109 ?
                      reg111 : {((reg113 ?
                              wire100 : reg107) * (reg115 >>> wire101)),
                          wire97})};
            end
          else
            begin
              reg119 <= {$signed(((&(|reg116)) >= {wire101}))};
              reg120 <= ($signed($unsigned($signed((wire100 ^~ wire98)))) ?
                  (($signed({reg116,
                      reg107}) <= $signed($unsigned(reg114))) ^~ (reg113 ?
                      reg113 : reg103[(1'h0):(1'h0)])) : ((($unsigned(reg104) ?
                          reg119 : reg120[(2'h3):(2'h2)]) - $signed((wire98 ?
                          wire101 : reg119))) ?
                      reg117[(3'h6):(3'h4)] : ($unsigned((-reg116)) << $signed((reg109 | reg116)))));
              reg121 <= $unsigned($signed(({(8'ha0)} ?
                  wire97 : (+$signed(wire97)))));
              reg122 <= ((((wire98 ^ (^~reg113)) ^~ $unsigned(reg113)) == {$unsigned($unsigned(reg117)),
                  (^~{reg106})}) | reg119[(1'h0):(1'h0)]);
              reg123 <= reg110;
            end
          reg124 <= reg118;
        end
    end
  assign wire125 = ((~^(-({(8'ha7)} ?
                       {(8'ha7)} : wire99))) < {$unsigned($signed({reg106,
                           wire98}))});
  assign wire126 = reg124[(3'h4):(3'h4)];
  always
    @(posedge clk) begin
      reg127 <= reg108[(2'h3):(1'h1)];
      if ($signed(reg104[(3'h5):(1'h0)]))
        begin
          reg128 <= {$signed($signed(($signed(reg122) >> ((8'hbe) ?
                  reg115 : reg109)))),
              (((-((8'hbc) && reg108)) ^~ (&reg121[(2'h3):(2'h3)])) ?
                  reg121 : $signed((wire100[(1'h0):(1'h0)] != reg119)))};
          if ((((8'hab) * $unsigned(reg113)) - $signed(((!$signed(wire100)) <= (wire99 ~^ (reg107 <= reg118))))))
            begin
              reg129 <= ((~|reg119) != $unsigned((reg107 ?
                  (reg128[(2'h2):(2'h2)] ?
                      (wire100 > wire101) : (~|reg124)) : ($signed(reg122) ?
                      (wire125 << (8'hba)) : (wire100 ? (8'had) : reg119)))));
              reg130 <= (7'h44);
              reg131 <= (!wire97);
            end
          else
            begin
              reg129 <= (8'hab);
              reg130 <= wire100;
              reg131 <= $signed((8'hbe));
            end
          reg132 <= ($unsigned(reg130) ?
              ($signed(($unsigned(reg120) ?
                  $unsigned(reg118) : $signed(reg108))) >= (wire101 ?
                  $unsigned(reg107) : $unsigned($signed(wire125)))) : (~(&wire97)));
          if (((reg117 >>> ((reg106 <= (reg113 ?
              reg111 : wire101)) <= reg115)) ^~ wire125))
            begin
              reg133 <= reg120[(4'hb):(2'h3)];
            end
          else
            begin
              reg133 <= (reg111[(3'h7):(1'h1)] ?
                  $signed(reg103[(4'h9):(3'h4)]) : $signed($unsigned($signed($unsigned(wire99)))));
              reg134 <= $signed(reg112);
              reg135 <= reg113[(3'h4):(1'h0)];
            end
        end
      else
        begin
          reg128 <= {$signed($signed(reg106)),
              $signed($unsigned((~|reg123[(2'h3):(2'h3)])))};
        end
    end
  assign wire136 = ((7'h44) ?
                       {(~$signed((reg115 ? reg111 : (8'hb4)))),
                           (|reg118)} : ({{$unsigned(reg102)}} <= reg127[(1'h1):(1'h1)]));
  assign wire137 = ({$unsigned(reg134)} ?
                       (8'ha5) : $unsigned($signed($unsigned((8'ha5)))));
  always
    @(posedge clk) begin
      reg138 <= wire96[(4'hf):(1'h1)];
      reg139 <= reg134;
      reg140 <= reg130[(1'h1):(1'h1)];
      reg141 <= reg129[(3'h6):(3'h5)];
      reg142 <= {reg113[(2'h2):(1'h1)]};
    end
  assign wire143 = (~|$signed((reg123[(3'h5):(1'h0)] ?
                       ((reg114 << reg130) >= (!reg120)) : reg102)));
  always
    @(posedge clk) begin
      if ((~|wire98))
        begin
          if ($unsigned(wire97[(1'h1):(1'h0)]))
            begin
              reg144 <= (((^~$signed((reg134 <<< wire125))) ?
                      (reg133 < (((8'haa) ? (8'ha0) : reg119) ?
                          reg104[(1'h0):(1'h0)] : $unsigned(reg114))) : $signed(reg108)) ?
                  (($signed($signed(wire98)) ?
                      {reg113[(4'h9):(3'h5)]} : reg102[(3'h6):(2'h3)]) + ({(wire125 ?
                              reg122 : reg130)} ?
                      reg115 : reg121)) : ((~&reg142) << reg104[(3'h5):(1'h1)]));
            end
          else
            begin
              reg144 <= $unsigned(reg133[(2'h2):(2'h2)]);
              reg145 <= $signed((&(+$signed(reg128[(3'h5):(1'h1)]))));
              reg146 <= reg128[(3'h4):(1'h0)];
            end
        end
      else
        begin
          reg144 <= reg140;
          reg145 <= (wire97 >> reg108);
          reg146 <= {$unsigned($signed((8'ha6)))};
          reg147 <= ($unsigned($signed(reg106[(3'h4):(1'h0)])) ?
              $signed(((reg118[(1'h0):(1'h0)] ?
                      (reg130 - reg145) : $signed(wire125)) ?
                  ((~&reg141) ?
                      ((8'hb8) ? reg124 : reg129) : (wire101 ?
                          (7'h42) : reg112)) : $unsigned({reg113,
                      (8'hb6)}))) : (~|$signed($unsigned((-(8'ha2))))));
        end
      reg148 <= (~|$signed((((8'hb0) ?
          (reg103 > (8'hb4)) : $unsigned(reg104)) >> reg110)));
      if (reg113)
        begin
          reg149 <= (^$unsigned((&$unsigned((reg119 >> reg141)))));
          if (reg111)
            begin
              reg150 <= $unsigned($signed(reg117));
              reg151 <= ({$unsigned($unsigned((wire125 ? reg119 : reg109)))} ?
                  {reg109[(4'ha):(4'h9)], (~|$signed({wire100}))} : reg108);
              reg152 <= $signed((|(^($unsigned(wire143) ?
                  $signed(reg119) : (&reg108)))));
              reg153 <= ($signed($signed($signed(reg146[(4'hc):(4'h9)]))) & {reg120[(4'hb):(1'h0)],
                  reg119});
              reg154 <= reg139[(2'h2):(2'h2)];
            end
          else
            begin
              reg150 <= {reg119[(3'h4):(1'h0)],
                  $unsigned((!($unsigned(wire99) ?
                      $unsigned(reg114) : {reg108, reg110})))};
              reg151 <= reg102;
              reg152 <= $unsigned(((((reg102 == reg121) ?
                      {reg123, reg146} : reg147[(4'ha):(4'ha)]) ?
                  (!reg144[(4'h9):(4'h8)]) : reg149[(1'h1):(1'h0)]) != $signed((~&reg108))));
              reg153 <= reg110;
              reg154 <= $signed(reg124[(4'hf):(4'hc)]);
            end
          reg155 <= (&$unsigned((((-(8'hb4)) ? $unsigned(reg112) : (+reg103)) ?
              reg131[(4'h8):(3'h4)] : $signed((&wire99)))));
          if ({($unsigned((8'ha2)) ? reg132 : {reg104})})
            begin
              reg156 <= reg124;
            end
          else
            begin
              reg156 <= ((+((reg123 ?
                  reg147 : $signed(reg150)) <= reg149[(3'h7):(1'h0)])) != $signed(reg110[(3'h4):(2'h2)]));
              reg157 <= (~|reg131);
              reg158 <= $unsigned($signed((reg155[(1'h0):(1'h0)] ?
                  $unsigned($unsigned(reg113)) : (reg142 && ((8'h9e) > wire96)))));
            end
        end
      else
        begin
          reg149 <= $unsigned($unsigned(reg138[(5'h14):(2'h2)]));
          reg150 <= (($signed($unsigned((&reg109))) ^ (~((reg132 ?
              reg109 : reg141) * reg105))) <= (+(+((^reg154) == $unsigned(reg105)))));
          reg151 <= $signed(($signed($signed($signed(reg107))) ?
              $signed(((wire126 | wire126) ?
                  reg138[(4'h9):(3'h6)] : ((8'hbd) ?
                      reg138 : (8'hbf)))) : reg158[(3'h6):(1'h0)]));
          if ((~(^($signed((reg107 ? reg149 : reg117)) ?
              (+(~&reg151)) : reg152))))
            begin
              reg152 <= ({($signed(reg116[(3'h7):(3'h4)]) ?
                      wire126 : (~{reg142})),
                  $signed($signed({reg145}))} >>> $unsigned(reg111));
              reg153 <= $unsigned(reg156);
              reg154 <= wire143;
              reg155 <= (({$signed($signed(reg114))} ~^ reg134) - (~$signed((reg119 ?
                  $signed(wire101) : (|reg153)))));
              reg156 <= reg119;
            end
          else
            begin
              reg152 <= (-$unsigned(reg116[(4'h8):(4'h8)]));
              reg153 <= ($unsigned($unsigned(reg146)) ?
                  (($signed(((8'ha5) <<< reg157)) ?
                      (reg127[(2'h3):(2'h3)] ?
                          (wire101 ?
                              reg135 : reg157) : $unsigned(reg127)) : ({reg120} ?
                          reg149 : ((8'hb2) ?
                              reg138 : wire97))) || ((-reg144[(4'h9):(3'h4)]) == reg130)) : (!($unsigned(reg111) ~^ {{(8'hb2),
                          (8'ha4)}})));
              reg154 <= (^~(reg151 ?
                  $unsigned({(reg147 <<< (8'ha7))}) : ($signed((8'hac)) || ($unsigned(reg148) || reg114[(1'h0):(1'h0)]))));
              reg155 <= $unsigned($signed(wire126[(3'h6):(2'h2)]));
            end
        end
      if ($signed(reg114[(1'h0):(1'h0)]))
        begin
          reg159 <= ((-(((reg133 ?
              (8'hb9) : wire99) ^~ $signed(reg102)) >> $signed($unsigned(reg114)))) < {{{$unsigned(reg107)},
                  $unsigned($unsigned(reg147))}});
          reg160 <= $unsigned((~reg145));
        end
      else
        begin
          if (({(8'hb3), reg142} & reg117[(3'h5):(2'h2)]))
            begin
              reg159 <= {$signed(reg115), wire125};
              reg160 <= {(!$signed($unsigned($signed(reg154))))};
              reg161 <= $signed({((+{(8'haa), reg123}) ?
                      ((wire99 + (8'hbf)) ?
                          (reg114 << reg127) : (8'ha6)) : $unsigned(reg112[(3'h7):(3'h6)]))});
              reg162 <= $signed($unsigned((((8'ha9) ?
                      {reg113, reg131} : (~reg146)) ?
                  $signed($signed(reg132)) : $signed({(8'hb9), reg146}))));
              reg163 <= reg117[(1'h0):(1'h0)];
            end
          else
            begin
              reg159 <= $signed($signed((wire101[(1'h1):(1'h1)] & $signed($signed(reg161)))));
              reg160 <= ($unsigned({$unsigned((reg113 ? reg134 : reg105)),
                  reg120[(4'hd):(4'hc)]}) | ($signed((7'h44)) <= {(reg115 <= reg133[(1'h1):(1'h0)]),
                  (reg140 ? $unsigned(reg111) : (reg121 ? wire100 : reg107))}));
              reg161 <= (8'hbe);
            end
          reg164 <= (-(reg117 >> reg138));
          reg165 <= reg149[(3'h5):(2'h3)];
        end
    end
  always
    @(posedge clk) begin
      reg166 <= ((+(+reg117[(3'h6):(2'h2)])) >= $unsigned((8'hac)));
      if (reg134)
        begin
          reg167 <= reg109;
          reg168 <= $unsigned($signed((((reg124 ?
              reg160 : reg113) << (reg129 + reg106)) <<< reg147[(4'hc):(2'h3)])));
          reg169 <= (reg166 | wire101);
        end
      else
        begin
          reg167 <= $unsigned((reg122 < $unsigned(($signed(reg148) <= (reg134 ~^ reg139)))));
          reg168 <= reg139;
          reg169 <= reg106;
          reg170 <= $unsigned($signed($unsigned(({(8'hac),
              reg145} | $signed(reg119)))));
        end
      reg171 <= $signed(reg108);
    end
  always
    @(posedge clk) begin
      reg172 <= $signed({{$signed((~|reg130)),
              {reg147[(5'h12):(3'h7)], (^(8'hb2))}},
          $unsigned($signed((reg132 & reg110)))});
    end
endmodule