(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param819 = (8'hb7))
(y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h1bf):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire4;
  input wire [(5'h10):(1'h0)] wire3;
  input wire [(5'h10):(1'h0)] wire2;
  input wire signed [(2'h3):(1'h0)] wire1;
  input wire [(3'h4):(1'h0)] wire0;
  wire [(3'h5):(1'h0)] wire818;
  reg [(4'hc):(1'h0)] reg817 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg816 = (1'h0);
  reg [(3'h7):(1'h0)] reg815 = (1'h0);
  reg [(4'h8):(1'h0)] reg814 = (1'h0);
  reg [(3'h7):(1'h0)] reg813 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg812 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg811 = (1'h0);
  reg [(5'h12):(1'h0)] forvar810 = (1'h0);
  reg [(5'h14):(1'h0)] reg809 = (1'h0);
  reg [(2'h2):(1'h0)] reg808 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg807 = (1'h0);
  reg [(4'h9):(1'h0)] reg806 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg805 = (1'h0);
  reg [(3'h4):(1'h0)] forvar804 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire802;
  wire signed [(4'hf):(1'h0)] wire628;
  wire signed [(4'hb):(1'h0)] wire28;
  reg signed [(3'h4):(1'h0)] reg27 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg26 = (1'h0);
  reg [(2'h3):(1'h0)] reg25 = (1'h0);
  reg [(4'hb):(1'h0)] reg24 = (1'h0);
  reg [(4'h9):(1'h0)] reg23 = (1'h0);
  reg [(2'h3):(1'h0)] reg22 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg21 = (1'h0);
  reg [(5'h12):(1'h0)] reg20 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar19 = (1'h0);
  reg [(5'h13):(1'h0)] reg18 = (1'h0);
  reg [(4'he):(1'h0)] reg17 = (1'h0);
  reg [(5'h12):(1'h0)] reg16 = (1'h0);
  reg [(3'h4):(1'h0)] reg15 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg14 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar13 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg12 = (1'h0);
  wire [(5'h15):(1'h0)] wire11;
  reg signed [(3'h6):(1'h0)] reg10 = (1'h0);
  reg [(5'h14):(1'h0)] reg9 = (1'h0);
  reg [(2'h3):(1'h0)] reg8 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg7 = (1'h0);
  reg [(5'h11):(1'h0)] reg6 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5 = (1'h0);
  assign y = {wire818,
                 reg817,
                 reg816,
                 reg815,
                 reg814,
                 reg813,
                 reg812,
                 reg811,
                 forvar810,
                 reg809,
                 reg808,
                 reg807,
                 reg806,
                 reg805,
                 forvar804,
                 wire802,
                 wire628,
                 wire28,
                 reg27,
                 reg26,
                 reg25,
                 reg24,
                 reg23,
                 reg22,
                 reg21,
                 reg20,
                 forvar19,
                 reg18,
                 reg17,
                 reg16,
                 reg15,
                 reg14,
                 forvar13,
                 reg12,
                 wire11,
                 reg10,
                 reg9,
                 reg8,
                 reg7,
                 reg6,
                 reg5,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg5 <= $unsigned(wire4[(3'h6):(3'h6)]);
      reg6 <= ((-$signed(wire0[(1'h1):(1'h0)])) >= wire3);
    end
  always
    @(posedge clk) begin
      reg7 <= wire1;
      reg8 <= (reg7[(4'hd):(4'hd)] ?
          $unsigned($signed(reg7[(3'h7):(2'h3)])) : {(8'hbc),
              reg7[(4'ha):(1'h1)]});
      reg9 <= (^~$unsigned((~^wire3)));
      reg10 = $unsigned((reg7 ? {wire4[(1'h1):(1'h0)], reg6} : reg9));
    end
  assign wire11 = {reg6};
  always
    @(posedge clk) begin
      reg12 = wire4;
      for (forvar13 = (1'h0); (forvar13 < (1'h0)); forvar13 = (forvar13 + (1'h1)))
        begin
          reg14 = (wire3[(3'h6):(3'h6)] <= reg5);
        end
    end
  always
    @(posedge clk) begin
      reg15 <= ((^~(($signed(reg12) ?
              (wire11 + reg10) : (-reg8)) ^ reg10[(1'h0):(1'h0)])) ?
          (wire3 ?
              $signed((!(wire11 ? reg6 : (8'ha9)))) : (wire4[(1'h0):(1'h0)] ?
                  (^~reg9[(4'hc):(2'h2)]) : {wire1, reg9})) : $unsigned(reg9));
    end
  always
    @(posedge clk) begin
      reg16 <= reg12[(4'he):(4'hc)];
      reg17 <= wire11[(4'h9):(2'h2)];
      reg18 <= $signed((|$signed($unsigned(reg15))));
    end
  always
    @(posedge clk) begin
      for (forvar19 = (1'h0); (forvar19 < (1'h0)); forvar19 = (forvar19 + (1'h1)))
        begin
          reg20 <= $unsigned($signed(reg16));
        end
      reg21 <= (8'hb8);
      reg22 = reg8;
      reg23 = (~&reg15[(1'h0):(1'h0)]);
      reg24 = (+$unsigned((8'h9d)));
    end
  always
    @(posedge clk) begin
      reg25 = ($unsigned($unsigned($unsigned($unsigned(reg10)))) >>> $signed({(^~(reg14 <<< reg12))}));
      reg26 <= ((^$unsigned($signed(reg14))) ?
          ($unsigned(((reg24 != forvar19) ?
              {(8'ha3), (8'ha2)} : forvar19)) | (($unsigned(reg22) ?
              $signed(reg7) : reg24) + reg23[(3'h5):(2'h2)])) : (&(+{(8'hb3)})));
      reg27 <= (forvar13[(1'h0):(1'h0)] ?
          reg7 : ($unsigned($unsigned(reg10)) && (~^reg20[(4'h8):(3'h7)])));
    end
  assign wire28 = $signed(reg8);
  module29 modinst629 (wire628, clk, wire4, reg21, reg6, reg24);
  module630 modinst803 (.y(wire802), .wire634(reg16), .wire632(wire628), .clk(clk), .wire631(wire28), .wire633(wire4));
  always
    @(posedge clk) begin
      for (forvar804 = (1'h0); (forvar804 < (1'h1)); forvar804 = (forvar804 + (1'h1)))
        begin
          reg805 = $unsigned({$unsigned(((8'ha7) ?
                  (wire1 ? reg22 : reg27) : $unsigned(reg7)))});
          reg806 <= ($unsigned(reg14) > ($signed(reg20[(3'h7):(2'h2)]) >= (~reg5[(3'h7):(3'h4)])));
          reg807 <= reg23[(4'h9):(4'h8)];
          reg808 <= ($signed(((+((7'h41) ? forvar804 : reg8)) <= (+reg21))) ?
              $signed($unsigned($unsigned((reg24 <<< reg21)))) : reg22);
        end
      reg809 <= (~reg14[(4'h8):(1'h0)]);
      for (forvar810 = (1'h0); (forvar810 < (1'h0)); forvar810 = (forvar810 + (1'h1)))
        begin
          if (({wire1} || {reg18}))
            begin
              reg811 <= reg12[(4'h8):(1'h0)];
              reg812 = $unsigned($unsigned(forvar13));
            end
          else
            begin
              reg811 <= {reg807,
                  $unsigned(($signed($signed(reg808)) == (!$unsigned(reg8))))};
              reg812 <= (((^~$unsigned(((8'ha6) ^~ reg18))) ?
                      (^~reg808) : forvar804[(1'h1):(1'h0)]) ?
                  (+reg21) : (wire11[(2'h2):(2'h2)] >> $signed({$signed(reg12),
                      $unsigned((8'hbc))})));
              reg813 <= (~$unsigned(reg25[(1'h0):(1'h0)]));
              reg814 <= reg16;
            end
          reg815 = $signed({{$signed((reg808 ? reg21 : reg15))}});
          reg816 <= reg5;
        end
      reg817 <= {($signed({$unsigned(forvar13), {reg808}}) ?
              reg17[(1'h0):(1'h0)] : ($signed((~^reg14)) ^~ $unsigned(wire628)))};
    end
  assign wire818 = reg20;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module630  (y, clk, wire631, wire632, wire633, wire634);
  output wire [(32'ha2):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hb):(1'h0)] wire631;
  input wire [(4'hf):(1'h0)] wire632;
  input wire signed [(5'h14):(1'h0)] wire633;
  input wire [(5'h12):(1'h0)] wire634;
  reg signed [(4'hc):(1'h0)] reg635 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg636 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg637 = (1'h0);
  reg [(3'h4):(1'h0)] reg638 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg639 = (1'h0);
  reg [(5'h13):(1'h0)] reg640 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg641 = (1'h0);
  wire [(4'h8):(1'h0)] wire642;
  reg [(5'h15):(1'h0)] reg643 = (1'h0);
  reg [(4'hb):(1'h0)] reg644 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg645 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire646;
  wire [(4'hd):(1'h0)] wire800;
  assign y = {reg635,
                 reg636,
                 reg637,
                 reg638,
                 reg639,
                 reg640,
                 reg641,
                 wire642,
                 reg643,
                 reg644,
                 reg645,
                 wire646,
                 wire800,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg635 <= $signed((^~wire633));
      if ($unsigned(((~|((8'hb9) != (|wire633))) ?
          {wire632[(4'h8):(4'h8)], (~wire634)} : ((&(wire631 ?
                  reg635 : reg635)) ?
              $signed((reg635 ?
                  wire634 : reg635)) : ((8'ha7) ^ ((8'ha8) & wire631))))))
        begin
          reg636 <= wire631[(3'h5):(1'h0)];
          reg637 <= $unsigned(($unsigned(wire634) - $signed(wire632[(4'h8):(2'h2)])));
          reg638 <= (^~((~(8'h9f)) || $unsigned($signed((reg637 ?
              reg636 : wire632)))));
        end
      else
        begin
          reg636 <= $signed($signed($unsigned(reg638[(1'h1):(1'h0)])));
          reg637 <= reg637;
          reg638 <= reg637[(4'ha):(4'h9)];
          reg639 <= wire632;
        end
      reg640 <= reg639[(1'h1):(1'h1)];
      reg641 <= (reg636[(2'h2):(1'h1)] ?
          $signed((reg637[(3'h5):(2'h3)] != wire634[(3'h6):(3'h4)])) : $signed((($signed(wire633) <= (reg640 != (7'h44))) >>> ((~^wire631) ?
              (reg635 ? (8'hbe) : (8'ha6)) : (+reg637)))));
    end
  assign wire642 = (8'had);
  always
    @(posedge clk) begin
      reg643 <= $unsigned({(~|($unsigned(reg636) - (-reg640)))});
      reg644 <= $signed((reg636[(4'hb):(4'h8)] ?
          (reg641[(3'h7):(3'h6)] && (+(reg638 <= reg640))) : ($unsigned($unsigned(reg638)) >= reg638)));
    end
  always
    @(posedge clk) begin
      reg645 <= (~^$signed(((~^((8'h9e) ? (8'h9d) : reg641)) ?
          reg635 : reg637[(4'hb):(3'h7)])));
    end
  assign wire646 = $signed((({wire633} ?
                       wire632 : $unsigned(wire633)) && ($signed((reg643 ^ wire631)) ?
                       ((~|reg636) && $signed(wire632)) : $signed({(8'hae),
                           wire634}))));
  module647 modinst801 (wire800, clk, reg643, reg640, wire634, reg635, reg644);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module29
#( parameter param626 = (^~(((+((8'hae) ? (8'ha6) : (8'haa))) ^ (((8'ha1) >> (8'ha8)) ? (|(7'h44)) : ((7'h44) ? (8'h9e) : (8'hbf)))) ? (8'hae) : (~&(((8'ha7) <<< (7'h42)) ? ((8'h9e) | (7'h44)) : (~|(8'had))))))
, parameter param627 = ((param626 || ({(~param626), (param626 ~^ param626)} ? ((param626 == param626) & (&(8'hba))) : ({param626} ? (param626 ? param626 : param626) : (8'hae)))) << {(param626 <= ((param626 ^ param626) ? (&param626) : (param626 ? param626 : (8'h9f)))), param626}) )
(y, clk, wire30, wire31, wire32, wire33);
  output wire [(32'h225):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire30;
  input wire signed [(4'h9):(1'h0)] wire31;
  input wire [(5'h11):(1'h0)] wire32;
  input wire [(4'hb):(1'h0)] wire33;
  wire signed [(5'h15):(1'h0)] wire34;
  reg signed [(2'h3):(1'h0)] forvar35 = (1'h0);
  reg [(5'h13):(1'h0)] reg36 = (1'h0);
  reg [(3'h7):(1'h0)] reg37 = (1'h0);
  reg [(5'h10):(1'h0)] reg38 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg39 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg40 = (1'h0);
  reg [(5'h10):(1'h0)] reg41 = (1'h0);
  reg [(4'he):(1'h0)] reg42 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg43 = (1'h0);
  reg [(4'hf):(1'h0)] forvar44 = (1'h0);
  reg [(3'h6):(1'h0)] reg45 = (1'h0);
  reg [(5'h15):(1'h0)] reg46 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire47;
  reg [(5'h13):(1'h0)] reg48 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg49 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg50 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg51 = (1'h0);
  reg [(3'h6):(1'h0)] forvar52 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar53 = (1'h0);
  reg [(3'h5):(1'h0)] reg54 = (1'h0);
  reg [(4'he):(1'h0)] reg55 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg56 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg57 = (1'h0);
  reg [(3'h4):(1'h0)] reg58 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg59 = (1'h0);
  reg [(4'hd):(1'h0)] forvar60 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg61 = (1'h0);
  reg [(2'h2):(1'h0)] reg62 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg63 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg64 = (1'h0);
  reg [(4'hf):(1'h0)] reg65 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg66 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg67 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg68 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg69 = (1'h0);
  reg [(5'h15):(1'h0)] reg70 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar65 = (1'h0);
  reg [(4'hd):(1'h0)] forvar71 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg72 = (1'h0);
  reg [(2'h3):(1'h0)] reg73 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar74 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg75 = (1'h0);
  reg [(5'h12):(1'h0)] reg76 = (1'h0);
  reg [(3'h7):(1'h0)] reg77 = (1'h0);
  wire [(4'ha):(1'h0)] wire368;
  wire [(4'ha):(1'h0)] wire370;
  wire [(2'h3):(1'h0)] wire624;
  assign y = {wire34,
                 forvar35,
                 reg36,
                 reg37,
                 reg38,
                 reg39,
                 reg40,
                 reg41,
                 reg42,
                 reg43,
                 forvar44,
                 reg45,
                 reg46,
                 wire47,
                 reg48,
                 reg49,
                 reg50,
                 reg51,
                 forvar52,
                 forvar53,
                 reg54,
                 reg55,
                 reg56,
                 reg57,
                 reg58,
                 reg59,
                 forvar60,
                 reg61,
                 reg62,
                 reg63,
                 reg64,
                 reg65,
                 reg66,
                 reg67,
                 reg68,
                 reg69,
                 reg70,
                 forvar65,
                 forvar71,
                 reg72,
                 reg73,
                 forvar74,
                 reg75,
                 reg76,
                 reg77,
                 wire368,
                 wire370,
                 wire624,
                 (1'h0)};
  assign wire34 = wire31;
  always
    @(posedge clk) begin
      for (forvar35 = (1'h0); (forvar35 < (1'h0)); forvar35 = (forvar35 + (1'h1)))
        begin
          reg36 <= {(~^wire33), (~|wire34[(4'hd):(4'hd)])};
          reg37 <= wire31[(3'h4):(1'h0)];
          reg38 <= wire32[(4'ha):(4'h8)];
          reg39 <= (~{(~$unsigned($signed(reg37))),
              (wire31[(1'h0):(1'h0)] ?
                  $unsigned({(8'ha7), reg37}) : $signed($signed(forvar35)))});
        end
      reg40 <= reg37[(3'h5):(1'h0)];
      reg41 <= reg39;
      reg42 <= {$unsigned(forvar35[(1'h1):(1'h0)])};
    end
  always
    @(posedge clk) begin
      reg43 <= $signed((&(7'h42)));
      for (forvar44 = (1'h0); (forvar44 < (1'h1)); forvar44 = (forvar44 + (1'h1)))
        begin
          reg45 <= (wire34 ?
              (8'ha9) : $unsigned((reg38 ?
                  reg37 : {reg42[(3'h7):(2'h2)], wire34})));
        end
      reg46 <= ($signed(((reg40 <<< {forvar44}) >> $unsigned((-wire33)))) ?
          reg41[(3'h5):(3'h5)] : reg39[(2'h2):(1'h0)]);
    end
  assign wire47 = ($unsigned(((reg40 ? wire34 : $unsigned(reg45)) ?
                          (~^(|reg46)) : $signed($signed(wire31)))) ?
                      $signed($unsigned(wire34[(3'h5):(1'h0)])) : $signed((reg37 ?
                          $unsigned({wire32, reg38}) : (((8'h9e) ?
                                  reg38 : reg39) ?
                              (reg41 ? (8'hb9) : wire31) : (-reg41)))));
  always
    @(posedge clk) begin
      reg48 <= $unsigned((reg43 ^~ $signed(((wire33 ? wire47 : reg38) - {reg38,
          forvar35}))));
      reg49 <= $signed(reg45[(1'h0):(1'h0)]);
      reg50 <= {reg43,
          (reg48 ?
              (|(((8'haf) | (8'hbc)) <= (wire34 <<< wire32))) : $signed($signed($signed(reg37))))};
      reg51 <= {(-reg45[(3'h4):(2'h3)]),
          {(&wire47), $signed($unsigned((wire33 ? reg42 : wire31)))}};
    end
  always
    @(posedge clk) begin
      for (forvar52 = (1'h0); (forvar52 < (1'h0)); forvar52 = (forvar52 + (1'h1)))
        begin
          for (forvar53 = (1'h0); (forvar53 < (3'h4)); forvar53 = (forvar53 + (1'h1)))
            begin
              reg54 <= reg48;
              reg55 <= reg50[(4'hc):(2'h2)];
            end
          reg56 = $signed(reg36[(2'h3):(1'h0)]);
        end
      reg57 <= {(($signed($unsigned((8'hbd))) == $unsigned($signed(reg36))) ?
              (($unsigned(forvar53) ~^ reg45) ?
                  $signed($signed(reg40)) : $signed({reg36})) : $unsigned(reg51)),
          (({(reg55 ? reg45 : reg49)} != $unsigned((^~reg51))) >= {(-{forvar35,
                  reg42}),
              ((!forvar52) <= (reg40 ? reg55 : reg42))})};
      reg58 <= $signed(wire33[(4'h9):(4'h9)]);
      reg59 <= (wire34[(4'he):(3'h5)] ?
          (~|$signed(reg43[(2'h2):(1'h1)])) : (reg56[(4'hd):(4'h8)] != wire32));
      for (forvar60 = (1'h0); (forvar60 < (1'h1)); forvar60 = (forvar60 + (1'h1)))
        begin
          reg61 <= {(wire31 ?
                  ($unsigned($unsigned((8'h9e))) <<< {((8'h9d) ?
                          reg58 : forvar60),
                      (|reg57)}) : {(~|reg57[(1'h0):(1'h0)]),
                      $signed(reg42[(4'hc):(3'h6)])}),
              ((!(^{reg46})) && (7'h40))};
          reg62 <= $unsigned(($unsigned(forvar60[(4'h9):(1'h0)]) ^ forvar53[(2'h2):(1'h0)]));
          reg63 <= (|$signed(reg37[(1'h1):(1'h0)]));
        end
    end
  always
    @(posedge clk) begin
      if ($unsigned(((^(wire47[(4'he):(4'he)] ?
              {forvar60, reg48} : (reg55 ? wire34 : wire32))) ?
          {$unsigned($signed((7'h44))),
              $unsigned($signed((7'h41)))} : {(reg58[(2'h3):(2'h2)] ?
                  (&wire31) : $unsigned(reg46)),
              ((7'h41) ? reg50[(5'h12):(4'hd)] : reg58[(2'h3):(1'h0)])})))
        begin
          reg64 <= (|(~|reg40[(1'h0):(1'h0)]));
          if ((reg55 ?
              wire31[(2'h3):(1'h1)] : (((reg39[(3'h5):(1'h0)] ?
                      reg36[(4'h9):(3'h5)] : $unsigned(forvar35)) ?
                  wire32 : ($signed(reg55) * {reg49})) >>> reg40)))
            begin
              reg65 <= $unsigned({{reg59,
                      ((reg50 ? reg58 : reg64) && (reg50 ? reg48 : reg64))}});
              reg66 <= reg58[(2'h3):(1'h1)];
              reg67 <= (+{(((~&wire31) == $unsigned(wire33)) || (((8'hb8) ?
                          (8'hb4) : reg51) ?
                      (reg54 ? reg50 : reg42) : $unsigned(reg38)))});
              reg68 <= $unsigned($unsigned((&reg48[(2'h3):(1'h1)])));
              reg69 = $unsigned({(~^((reg45 ? reg48 : wire32) && (-(8'h9c))))});
            end
          else
            begin
              reg65 <= ($signed($unsigned(($unsigned(wire34) ?
                  reg40 : (reg38 >>> reg48)))) == reg45[(1'h1):(1'h1)]);
              reg66 <= $signed({((~&$signed(reg55)) ?
                      reg43[(2'h3):(1'h1)] : $unsigned((reg64 * reg49))),
                  ((~^(7'h41)) ?
                      $signed(reg45) : $unsigned((wire33 || reg61)))});
              reg67 = ((8'h9e) & $unsigned(reg59));
              reg68 <= $unsigned($unsigned((7'h44)));
              reg69 <= reg59[(1'h0):(1'h0)];
            end
          reg70 = $unsigned((8'h9d));
        end
      else
        begin
          reg64 <= (reg38 < (($unsigned((reg69 ?
              reg70 : reg46)) >>> ($signed(reg49) ?
              (wire32 > (8'ha4)) : (+reg67))) != $unsigned(reg66[(4'hf):(1'h0)])));
          for (forvar65 = (1'h0); (forvar65 < (2'h3)); forvar65 = (forvar65 + (1'h1)))
            begin
              reg66 <= {$unsigned((($signed(reg62) >>> reg70[(3'h7):(1'h0)]) ?
                      {$unsigned(reg38), {reg58}} : $unsigned(reg57))),
                  (reg43[(1'h0):(1'h0)] <<< (forvar35 != $signed((reg67 ?
                      wire33 : reg49))))};
              reg67 = ($signed(forvar52) ?
                  {(8'h9d),
                      ({reg64[(2'h3):(2'h3)]} ?
                          (!reg48) : (~&(~reg65)))} : reg37[(3'h5):(1'h1)]);
              reg68 <= reg69;
            end
          reg69 <= $signed(reg56);
        end
      for (forvar71 = (1'h0); (forvar71 < (1'h1)); forvar71 = (forvar71 + (1'h1)))
        begin
          reg72 <= (((((wire30 ? reg48 : reg41) ?
                      $unsigned(reg57) : $signed((8'hb1))) & reg68[(3'h7):(3'h4)]) ?
                  $signed((reg69 ^ reg55[(2'h2):(1'h0)])) : $unsigned({(8'hac),
                      $signed(reg51)})) ?
              (^~$unsigned(reg39)) : reg62[(1'h0):(1'h0)]);
          reg73 <= (reg66 ?
              $signed(($unsigned((reg62 ? (8'ha5) : (8'hbf))) ?
                  ((reg64 << forvar35) ?
                      reg57[(2'h3):(2'h3)] : (forvar71 >= reg42)) : ((reg58 ?
                          forvar44 : reg66) ?
                      $signed(reg67) : (reg72 ^ reg54)))) : {((&forvar52) ?
                      $signed($unsigned(reg62)) : $unsigned($signed(reg49)))});
          for (forvar74 = (1'h0); (forvar74 < (2'h3)); forvar74 = (forvar74 + (1'h1)))
            begin
              reg75 <= reg65[(4'hf):(4'he)];
              reg76 <= (~{$unsigned(({forvar74,
                      wire47} ~^ forvar71[(4'hc):(4'h8)])),
                  (8'hb1)});
              reg77 <= $unsigned({(&((^~reg45) && (reg68 & forvar52))),
                  reg48[(4'ha):(2'h3)]});
            end
        end
    end
  module78 modinst369 (wire368, clk, reg41, forvar65, reg70, forvar44);
  assign wire370 = {(~&forvar35),
                       ($signed((!(forvar74 == forvar71))) <= $unsigned((!$signed(reg37))))};
  module371 modinst625 (.wire372(reg65), .wire376(reg61), .wire375(reg77), .clk(clk), .y(wire624), .wire373(reg46), .wire374(reg40));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module371  (y, clk, wire376, wire375, wire374, wire373, wire372);
  output wire [(32'h39f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire376;
  input wire [(3'h7):(1'h0)] wire375;
  input wire [(4'ha):(1'h0)] wire374;
  input wire signed [(5'h15):(1'h0)] wire373;
  input wire [(4'hc):(1'h0)] wire372;
  reg signed [(2'h2):(1'h0)] reg623 = (1'h0);
  reg [(4'hb):(1'h0)] reg622 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg621 = (1'h0);
  reg [(4'hc):(1'h0)] forvar620 = (1'h0);
  reg [(4'hc):(1'h0)] reg619 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg618 = (1'h0);
  reg [(4'hc):(1'h0)] reg617 = (1'h0);
  reg [(3'h5):(1'h0)] reg616 = (1'h0);
  reg [(5'h15):(1'h0)] reg615 = (1'h0);
  reg [(3'h6):(1'h0)] reg614 = (1'h0);
  reg [(4'hd):(1'h0)] forvar613 = (1'h0);
  reg [(4'hd):(1'h0)] reg612 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar611 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg610 = (1'h0);
  wire [(4'hc):(1'h0)] wire609;
  wire signed [(5'h15):(1'h0)] wire608;
  wire signed [(3'h5):(1'h0)] wire607;
  wire signed [(4'ha):(1'h0)] wire606;
  reg signed [(5'h10):(1'h0)] reg605 = (1'h0);
  reg [(2'h2):(1'h0)] reg604 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg603 = (1'h0);
  reg [(4'hb):(1'h0)] reg602 = (1'h0);
  reg [(4'he):(1'h0)] reg601 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar600 = (1'h0);
  reg [(4'he):(1'h0)] reg599 = (1'h0);
  reg [(5'h13):(1'h0)] reg598 = (1'h0);
  reg [(2'h2):(1'h0)] reg597 = (1'h0);
  reg [(5'h12):(1'h0)] forvar596 = (1'h0);
  reg [(3'h7):(1'h0)] reg595 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg594 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg593 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg592 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar591 = (1'h0);
  reg [(4'ha):(1'h0)] reg590 = (1'h0);
  reg [(5'h15):(1'h0)] reg589 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire588;
  reg [(4'h8):(1'h0)] reg587 = (1'h0);
  reg [(3'h4):(1'h0)] reg586 = (1'h0);
  reg [(4'hf):(1'h0)] reg585 = (1'h0);
  reg [(2'h3):(1'h0)] reg584 = (1'h0);
  wire [(4'hd):(1'h0)] wire583;
  reg signed [(4'he):(1'h0)] reg582 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg581 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg580 = (1'h0);
  reg [(3'h5):(1'h0)] reg579 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg578 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg577 = (1'h0);
  reg [(4'hb):(1'h0)] reg576 = (1'h0);
  reg [(5'h14):(1'h0)] reg575 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg574 = (1'h0);
  reg [(4'hb):(1'h0)] reg573 = (1'h0);
  reg [(2'h2):(1'h0)] reg572 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg571 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg570 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar569 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg568 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg567 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar566 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg565 = (1'h0);
  reg [(2'h2):(1'h0)] reg564 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg563 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar562 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg561 = (1'h0);
  reg [(4'hf):(1'h0)] reg560 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar559 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg558 = (1'h0);
  reg [(4'he):(1'h0)] reg557 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg556 = (1'h0);
  reg [(4'hc):(1'h0)] reg555 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar554 = (1'h0);
  wire [(5'h14):(1'h0)] wire553;
  wire [(4'hc):(1'h0)] wire552;
  reg [(3'h4):(1'h0)] reg551 = (1'h0);
  reg [(3'h4):(1'h0)] reg550 = (1'h0);
  reg [(4'he):(1'h0)] forvar549 = (1'h0);
  reg [(2'h3):(1'h0)] reg548 = (1'h0);
  reg [(3'h6):(1'h0)] reg547 = (1'h0);
  reg [(4'ha):(1'h0)] reg546 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg545 = (1'h0);
  reg [(5'h11):(1'h0)] reg544 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg543 = (1'h0);
  reg [(5'h15):(1'h0)] reg542 = (1'h0);
  reg [(2'h2):(1'h0)] reg541 = (1'h0);
  wire [(3'h4):(1'h0)] wire539;
  assign y = {reg623,
                 reg622,
                 reg621,
                 forvar620,
                 reg619,
                 reg618,
                 reg617,
                 reg616,
                 reg615,
                 reg614,
                 forvar613,
                 reg612,
                 forvar611,
                 reg610,
                 wire609,
                 wire608,
                 wire607,
                 wire606,
                 reg605,
                 reg604,
                 reg603,
                 reg602,
                 reg601,
                 forvar600,
                 reg599,
                 reg598,
                 reg597,
                 forvar596,
                 reg595,
                 reg594,
                 reg593,
                 reg592,
                 forvar591,
                 reg590,
                 reg589,
                 wire588,
                 reg587,
                 reg586,
                 reg585,
                 reg584,
                 wire583,
                 reg582,
                 reg581,
                 reg580,
                 reg579,
                 reg578,
                 reg577,
                 reg576,
                 reg575,
                 reg574,
                 reg573,
                 reg572,
                 reg571,
                 reg570,
                 forvar569,
                 reg568,
                 reg567,
                 forvar566,
                 reg565,
                 reg564,
                 reg563,
                 forvar562,
                 reg561,
                 reg560,
                 forvar559,
                 reg558,
                 reg557,
                 reg556,
                 reg555,
                 forvar554,
                 wire553,
                 wire552,
                 reg551,
                 reg550,
                 forvar549,
                 reg548,
                 reg547,
                 reg546,
                 reg545,
                 reg544,
                 reg543,
                 reg542,
                 reg541,
                 wire539,
                 (1'h0)};
  module377 modinst540 (.wire378(wire373), .wire381(wire372), .wire380(wire376), .wire379(wire374), .clk(clk), .y(wire539));
  always
    @(posedge clk) begin
      reg541 = wire539;
    end
  always
    @(posedge clk) begin
      reg542 <= ($unsigned($signed((wire375[(2'h3):(1'h0)] ?
              wire372[(4'h9):(3'h6)] : (+wire539)))) ?
          $signed($signed(((wire375 << wire374) ?
              (^wire376) : wire373[(4'hb):(3'h5)]))) : (wire374[(4'ha):(4'h8)] ?
              (wire372 ^~ $signed((!wire373))) : (($unsigned(wire375) + (wire372 ^ wire373)) ?
                  wire373 : (|$unsigned(wire373)))));
      reg543 = wire373;
    end
  always
    @(posedge clk) begin
      reg544 <= wire374;
      reg545 <= reg544;
      reg546 <= (8'hb6);
      reg547 = {$unsigned($unsigned({$unsigned((8'haf)), $signed(reg541)})),
          {(reg545 ?
                  reg543[(3'h4):(2'h3)] : {(wire372 && reg545),
                      $unsigned((8'ha6))})}};
      reg548 <= (wire372 ~^ wire375);
    end
  always
    @(posedge clk) begin
      for (forvar549 = (1'h0); (forvar549 < (1'h0)); forvar549 = (forvar549 + (1'h1)))
        begin
          reg550 <= wire376[(4'hd):(4'hc)];
        end
      reg551 <= (8'hac);
    end
  assign wire552 = reg544;
  assign wire553 = (~^(!$unsigned($unsigned(reg551[(2'h2):(1'h0)]))));
  always
    @(posedge clk) begin
      for (forvar554 = (1'h0); (forvar554 < (1'h0)); forvar554 = (forvar554 + (1'h1)))
        begin
          reg555 <= reg542;
        end
      reg556 <= (|(~&(((+forvar549) ?
          wire539[(1'h0):(1'h0)] : ((8'h9d) ? reg545 : wire373)) != (8'h9f))));
      reg557 <= reg555;
      reg558 <= (8'hb9);
      for (forvar559 = (1'h0); (forvar559 < (2'h3)); forvar559 = (forvar559 + (1'h1)))
        begin
          reg560 = wire553;
          reg561 = (8'hb8);
          for (forvar562 = (1'h0); (forvar562 < (1'h0)); forvar562 = (forvar562 + (1'h1)))
            begin
              reg563 <= (reg556 < $signed($signed((7'h42))));
              reg564 <= (($signed(wire375) >>> reg558[(3'h5):(3'h5)]) <<< $signed(reg542));
              reg565 <= ($signed(reg555) ?
                  (((reg548[(2'h3):(2'h3)] != {(8'hbc)}) != (^(reg557 ?
                      wire373 : (8'ha2)))) | forvar562) : {reg547[(3'h4):(1'h0)],
                      (((8'hb1) && (!reg564)) == $unsigned(((8'hac) ?
                          reg555 : reg550)))});
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar566 = (1'h0); (forvar566 < (1'h0)); forvar566 = (forvar566 + (1'h1)))
        begin
          reg567 = {({$signed((wire553 * wire552))} - $signed($unsigned((wire374 + forvar554)))),
              (8'ha5)};
          reg568 <= reg567[(3'h4):(1'h0)];
          for (forvar569 = (1'h0); (forvar569 < (1'h1)); forvar569 = (forvar569 + (1'h1)))
            begin
              reg570 = $signed(({(~&wire539[(2'h3):(1'h0)])} >> forvar569[(1'h1):(1'h1)]));
              reg571 <= forvar566;
              reg572 <= $unsigned((!reg567[(3'h4):(2'h3)]));
            end
          reg573 <= (($unsigned($signed(wire372)) < $signed(((8'hb8) ~^ $signed((8'hb1))))) <= $unsigned({{$unsigned(forvar566)},
              ($signed(reg567) ^~ $unsigned(wire372))}));
        end
      reg574 <= (($signed((reg568 ? wire553 : wire539)) ?
          reg542[(5'h15):(4'hc)] : reg567) <<< $signed(wire372[(3'h7):(1'h0)]));
      reg575 = ($signed(($unsigned((~&forvar549)) ^~ $signed({reg541}))) >= reg573[(4'hb):(3'h6)]);
      reg576 <= reg544;
      reg577 <= (8'h9d);
    end
  always
    @(posedge clk) begin
      reg578 = (((((reg568 ?
              reg573 : reg560) << (&(8'hb8))) >> (~$signed((8'ha1)))) ~^ ({$signed((8'haf)),
              reg575} >>> $signed((wire375 ? forvar562 : wire374)))) ?
          reg573 : $signed($unsigned((~&{reg543, reg570}))));
      reg579 <= forvar549[(4'hb):(2'h2)];
      reg580 = $signed({wire539[(2'h2):(1'h1)],
          ({{reg578, reg568}} ? wire552 : (&$signed(reg547)))});
      reg581 <= forvar549;
      reg582 <= $unsigned({$signed(($signed(reg575) ?
              $unsigned(reg547) : wire372[(4'hb):(3'h4)])),
          reg573[(3'h5):(3'h5)]});
    end
  assign wire583 = (((~wire376) ?
                       (~|(forvar549 || (^~reg578))) : (forvar549[(4'ha):(1'h0)] ^~ reg577)) == $signed($signed(((reg577 & forvar569) ?
                       (reg574 ? reg551 : reg561) : (|reg564)))));
  always
    @(posedge clk) begin
      reg584 = ((^~(~($unsigned(reg546) ?
              reg551[(1'h1):(1'h1)] : $signed(reg555)))) ?
          wire374 : {((forvar559 ? reg581[(1'h1):(1'h0)] : {reg543, (8'hae)}) ?
                  ($signed(reg579) ?
                      (reg574 * reg551) : forvar566[(5'h11):(4'hd)]) : reg547),
              (&{(wire373 ? reg575 : (8'h9f)), {reg563}})});
      reg585 = (8'haf);
      reg586 <= $unsigned($signed(forvar549));
      reg587 <= reg557;
    end
  assign wire588 = ((^reg581) < {$unsigned($unsigned($unsigned(wire553))),
                       (~|$signed(wire553[(3'h5):(2'h3)]))});
  always
    @(posedge clk) begin
      reg589 <= reg542;
      reg590 <= {(((forvar566 ?
              (reg567 != reg567) : $unsigned(reg589)) <= ((reg544 >>> wire376) ?
              ((8'hb8) <<< reg580) : $unsigned(reg572))) * ($unsigned((~^reg580)) != reg565[(2'h2):(1'h1)]))};
      for (forvar591 = (1'h0); (forvar591 < (1'h1)); forvar591 = (forvar591 + (1'h1)))
        begin
          reg592 <= $signed($unsigned(reg580[(4'hc):(4'h8)]));
          reg593 <= ($unsigned(forvar591[(3'h6):(2'h2)]) ?
              $signed(reg574[(4'hb):(2'h3)]) : (|$unsigned($signed($unsigned(wire372)))));
          reg594 <= (~&reg573[(3'h5):(1'h0)]);
        end
      reg595 <= forvar554[(4'hd):(1'h0)];
      for (forvar596 = (1'h0); (forvar596 < (1'h1)); forvar596 = (forvar596 + (1'h1)))
        begin
          reg597 <= reg543[(1'h1):(1'h1)];
          reg598 <= reg568[(4'h8):(4'h8)];
          reg599 <= ((reg567[(2'h3):(2'h3)] ?
              $signed(reg579[(1'h0):(1'h0)]) : {(!{reg561}),
                  (-reg563[(3'h6):(3'h5)])}) << ((|forvar569[(3'h5):(1'h0)]) ?
              $signed(reg580) : {$unsigned((forvar562 ? wire583 : (7'h41)))}));
          for (forvar600 = (1'h0); (forvar600 < (2'h3)); forvar600 = (forvar600 + (1'h1)))
            begin
              reg601 <= (((8'hb5) ?
                  ($signed(reg577[(2'h3):(2'h3)]) + $unsigned((!(7'h42)))) : $unsigned(((reg593 ?
                          reg545 : reg541) ?
                      $unsigned(reg545) : wire376[(4'hf):(2'h3)]))) == ((~^{(|reg578),
                  ((8'hb1) ?
                      (8'ha0) : reg551)}) >= (~$unsigned($unsigned(reg567)))));
              reg602 <= ((forvar569[(1'h1):(1'h1)] ?
                  $unsigned((reg597[(1'h1):(1'h1)] && $signed(reg541))) : (((reg541 ?
                      (7'h44) : forvar600) <<< $unsigned(forvar549)) != $signed((+reg581)))) > ({wire376[(4'ha):(4'h8)]} ?
                  $signed($unsigned($signed((8'hb5)))) : ({(!reg556)} ?
                      ((+(8'haf)) + reg578) : ((|wire539) ?
                          $signed(reg584) : reg580))));
              reg603 <= (((((reg556 ^ reg564) ?
                          (^reg550) : reg557) ^~ $signed($signed(wire588))) ?
                      (~&{(reg587 ^~ reg550), (~^reg567)}) : (((reg593 ?
                              reg546 : (8'hbf)) || reg570[(3'h5):(1'h0)]) ?
                          ((^~reg585) ?
                              reg575[(5'h14):(2'h3)] : reg590[(1'h1):(1'h0)]) : ({reg573,
                                  reg595} ?
                              reg576[(2'h3):(1'h0)] : reg582[(4'ha):(2'h3)]))) ?
                  ((~^(~|(8'ha3))) ?
                      reg586[(1'h1):(1'h0)] : $unsigned((wire539[(2'h3):(1'h0)] >> (!wire553)))) : (8'hbc));
              reg604 <= (reg587 << (^(^($signed(reg601) > {reg592, wire373}))));
              reg605 = reg580[(4'h9):(3'h6)];
            end
        end
    end
  assign wire606 = (({(~|forvar566)} ?
                       (~((-wire539) ?
                           forvar591 : $unsigned(forvar596))) : wire372[(4'h8):(3'h7)]) != reg557);
  assign wire607 = reg555[(1'h1):(1'h1)];
  assign wire608 = ((~&wire376[(3'h6):(3'h5)]) ?
                       (((wire539[(1'h0):(1'h0)] ?
                                   $signed((8'hae)) : reg601[(4'hd):(3'h5)]) ?
                               $unsigned({reg593, (8'ha1)}) : (&(!reg560))) ?
                           $signed(reg545[(4'h8):(4'h8)]) : (reg602 > (~&$unsigned((8'ha5))))) : forvar596[(5'h11):(3'h4)]);
  assign wire609 = reg587;
  always
    @(posedge clk) begin
      reg610 <= wire609;
      for (forvar611 = (1'h0); (forvar611 < (3'h4)); forvar611 = (forvar611 + (1'h1)))
        begin
          reg612 <= reg604[(2'h2):(1'h0)];
          for (forvar613 = (1'h0); (forvar613 < (1'h1)); forvar613 = (forvar613 + (1'h1)))
            begin
              reg614 <= $unsigned($unsigned(reg612[(4'hc):(2'h2)]));
              reg615 <= ($signed({((-reg561) ?
                      $unsigned(reg586) : (reg576 ?
                          reg612 : (8'hbd)))}) - ($unsigned($unsigned($signed(reg585))) ?
                  $signed(((reg594 && wire608) * (reg574 ?
                      wire373 : reg598))) : {((reg561 > (8'h9d)) << reg546[(1'h1):(1'h1)])}));
              reg616 = reg543;
              reg617 <= (+$unsigned((^~$signed($unsigned(reg560)))));
            end
          reg618 = $signed(($signed((reg612[(3'h7):(2'h3)] ?
              (reg543 | reg567) : $signed((8'hba)))) >= ((|reg563[(4'h8):(3'h4)]) ?
              (wire553[(1'h0):(1'h0)] ?
                  $signed(forvar554) : (|wire552)) : wire373)));
        end
      reg619 = (~|(reg550[(3'h4):(3'h4)] ?
          (reg578 ^ $signed({reg612})) : reg574[(4'hc):(3'h4)]));
      for (forvar620 = (1'h0); (forvar620 < (3'h4)); forvar620 = (forvar620 + (1'h1)))
        begin
          reg621 <= $unsigned($unsigned((((forvar549 ^~ reg597) ?
              reg570[(2'h3):(1'h0)] : $signed(reg551)) || (7'h41))));
          reg622 <= wire552[(3'h6):(3'h5)];
        end
      reg623 = reg612;
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module78  (y, clk, wire82, wire81, wire80, wire79);
  output wire [(32'h18f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire82;
  input wire [(4'hf):(1'h0)] wire81;
  input wire [(4'h9):(1'h0)] wire80;
  input wire signed [(4'hf):(1'h0)] wire79;
  reg [(4'he):(1'h0)] reg367 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg366 = (1'h0);
  reg [(2'h2):(1'h0)] reg365 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg364 = (1'h0);
  reg [(4'hc):(1'h0)] reg363 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar362 = (1'h0);
  reg [(4'hf):(1'h0)] reg361 = (1'h0);
  reg [(4'h8):(1'h0)] forvar360 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg359 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg358 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg357 = (1'h0);
  reg [(4'hc):(1'h0)] reg356 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg355 = (1'h0);
  reg [(4'hd):(1'h0)] forvar354 = (1'h0);
  wire [(4'he):(1'h0)] wire353;
  wire [(4'hd):(1'h0)] wire352;
  wire signed [(5'h15):(1'h0)] wire350;
  reg [(5'h11):(1'h0)] reg284 = (1'h0);
  reg [(4'hf):(1'h0)] reg283 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg282 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg281 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire280;
  wire signed [(4'ha):(1'h0)] wire278;
  reg signed [(4'hd):(1'h0)] reg110 = (1'h0);
  reg [(4'hd):(1'h0)] reg109 = (1'h0);
  reg [(5'h13):(1'h0)] reg108 = (1'h0);
  reg [(2'h2):(1'h0)] reg107 = (1'h0);
  reg [(2'h3):(1'h0)] reg106 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg105 = (1'h0);
  reg [(5'h13):(1'h0)] reg104 = (1'h0);
  reg [(4'h9):(1'h0)] reg103 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire101;
  assign y = {reg367,
                 reg366,
                 reg365,
                 reg364,
                 reg363,
                 forvar362,
                 reg361,
                 forvar360,
                 reg359,
                 reg358,
                 reg357,
                 reg356,
                 reg355,
                 forvar354,
                 wire353,
                 wire352,
                 wire350,
                 reg284,
                 reg283,
                 reg282,
                 reg281,
                 wire280,
                 wire278,
                 reg110,
                 reg109,
                 reg108,
                 reg107,
                 reg106,
                 reg105,
                 reg104,
                 reg103,
                 wire101,
                 (1'h0)};
  module83 modinst102 (.wire85(wire82), .clk(clk), .wire86(wire81), .wire84((8'ha1)), .y(wire101), .wire87(wire79), .wire88(wire80));
  always
    @(posedge clk) begin
      reg103 = $unsigned((~$unsigned((|$signed(wire80)))));
      reg104 = $signed(wire101[(3'h5):(1'h0)]);
      reg105 <= (reg103 * $signed(wire79[(4'hc):(2'h3)]));
    end
  always
    @(posedge clk) begin
      reg106 <= $signed($unsigned((reg105 ?
          $unsigned(reg104) : ((8'hac) ? (wire80 & (8'h9f)) : (+(8'hb8))))));
      reg107 <= ($signed((-reg106)) + wire101);
      reg108 <= (wire101[(1'h1):(1'h1)] > (~^(-$unsigned((^~reg106)))));
      reg109 <= (^$unsigned($signed($unsigned((8'hb9)))));
      reg110 = (~|($unsigned(wire81) > $signed(reg105)));
    end
  module111 modinst279 (wire278, clk, reg105, reg104, reg108, reg109);
  assign wire280 = (reg105[(5'h12):(4'he)] < $unsigned($signed($signed((+reg110)))));
  always
    @(posedge clk) begin
      reg281 <= reg108[(4'h8):(1'h0)];
      reg282 <= (|reg104);
      reg283 <= reg109;
      reg284 <= (+({(~&$signed(reg103)), reg281} ?
          ($signed({reg108, (8'ha1)}) ?
              reg103[(3'h6):(1'h1)] : {(reg110 >> (8'hbe))}) : $unsigned($unsigned($signed(wire79)))));
    end
  module285 modinst351 (wire350, clk, wire81, wire280, wire101, reg109);
  assign wire352 = $unsigned({$unsigned(((reg104 <= reg281) ?
                           $unsigned(wire79) : $signed(reg282)))});
  assign wire353 = (wire352 < (reg105[(5'h13):(4'ha)] ?
                       $signed($unsigned($unsigned(reg110))) : (wire81[(2'h3):(2'h2)] ?
                           $unsigned(wire278) : ((~|wire350) >= (wire278 > wire352)))));
  always
    @(posedge clk) begin
      for (forvar354 = (1'h0); (forvar354 < (1'h1)); forvar354 = (forvar354 + (1'h1)))
        begin
          reg355 <= $signed(reg283);
          reg356 <= $signed((($unsigned({wire82,
                  reg283}) <<< $signed($signed(wire280))) ?
              ($unsigned($signed(reg281)) >= {$unsigned(wire352)}) : wire81));
          reg357 <= reg110[(2'h2):(1'h0)];
          reg358 = {{(($signed(reg281) ?
                      reg357[(1'h1):(1'h1)] : (^~reg104)) <<< ((!wire280) ?
                      reg106 : (wire101 ? reg284 : wire353))),
                  wire101[(4'hd):(4'h9)]}};
          reg359 = ($unsigned($unsigned(wire353)) ^ $signed(({((8'haf) ?
                  reg358 : reg281)} > $signed((reg357 <= reg107)))));
        end
      for (forvar360 = (1'h0); (forvar360 < (2'h3)); forvar360 = (forvar360 + (1'h1)))
        begin
          reg361 = ($unsigned((((reg104 ?
                  reg284 : wire82) >> $unsigned(reg357)) ?
              ($signed(reg110) ?
                  $signed((8'hae)) : $signed((8'hbf))) : (+((8'hbd) < forvar354)))) ^ ((~&{{(8'h9d)}}) & $signed($signed({forvar354}))));
        end
      for (forvar362 = (1'h0); (forvar362 < (1'h1)); forvar362 = (forvar362 + (1'h1)))
        begin
          reg363 = ({{$unsigned($signed(reg283)), (~&(~forvar362))}} ?
              wire82 : $signed((~^(|reg104[(4'he):(2'h3)]))));
          reg364 <= (~&$unsigned(wire80));
          reg365 <= ($signed((reg355 ?
                  (reg283 ? (+(8'ha5)) : $unsigned((8'had))) : (&{wire79}))) ?
              $signed({{reg361}}) : {($unsigned((-(8'hb2))) ?
                      reg364[(3'h6):(1'h1)] : $unsigned($unsigned(wire352)))});
        end
      reg366 <= ((^(reg110[(2'h3):(1'h0)] ?
              reg356[(3'h5):(3'h4)] : (-$signed(reg284)))) ?
          wire80[(1'h0):(1'h0)] : ((reg357[(1'h0):(1'h0)] ?
              (8'ha0) : reg105[(3'h4):(1'h1)]) > (({wire101} ^~ $signed(reg358)) ?
              reg361 : (+forvar362))));
      reg367 <= $unsigned(reg105);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module285
#( parameter param348 = (((({(8'hb9)} == (8'hb8)) <<< {{(8'h9c)}, {(8'hac), (8'hb0)}}) >> (({(8'h9c)} ? (~&(8'hae)) : ((8'ha0) ? (8'hbd) : (8'ha4))) ? (~&((8'had) < (8'hb2))) : (-(+(7'h43))))) ? (((((8'hb7) == (8'hb4)) ? ((8'ha7) > (8'ha8)) : {(8'hab)}) >= (((8'hb3) == (7'h43)) != ((8'hbc) == (8'ha7)))) ? {({(8'ha6)} ? (^~(7'h40)) : ((8'ha2) - (8'hb0))), ((^(8'hb5)) ^ (!(7'h42)))} : ((((8'hb9) ~^ (8'had)) * ((8'hae) ? (8'h9f) : (8'haa))) <<< ((^~(8'ha3)) ? {(8'ha6)} : ((8'ha2) != (8'hbf))))) : (((^{(8'haa), (8'ha4)}) ? (^(|(7'h41))) : (!((8'h9d) ? (8'hb2) : (8'hbc)))) ? (((+(7'h43)) ~^ (8'hba)) ? (~^(+(7'h43))) : ({(8'hb5)} == ((8'hbc) ? (8'hb1) : (8'hab)))) : (~^{((8'ha4) << (8'haf))})))
, parameter param349 = ((&{(~^(param348 ? (7'h41) : (8'ha3)))}) ? (((-(param348 >= param348)) ? ({param348, param348} ? {param348, param348} : ((8'hb9) ^~ param348)) : ((^param348) | param348)) ? {(~^(param348 || param348)), ((param348 ^~ param348) ? param348 : (~param348))} : (((param348 ? param348 : param348) ^~ (param348 ? param348 : param348)) - ({param348} <<< param348))) : {(param348 ? ((param348 ? param348 : param348) ? (8'ha5) : {param348, param348}) : param348), (^{(~&param348)})}) )
(y, clk, wire289, wire288, wire287, wire286);
  output wire [(32'h2d6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire289;
  input wire signed [(5'h11):(1'h0)] wire288;
  input wire signed [(5'h10):(1'h0)] wire287;
  input wire signed [(3'h6):(1'h0)] wire286;
  wire [(2'h2):(1'h0)] wire347;
  wire [(4'hd):(1'h0)] wire346;
  reg [(3'h6):(1'h0)] reg345 = (1'h0);
  reg [(4'hd):(1'h0)] reg344 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg343 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg342 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg341 = (1'h0);
  reg [(4'h8):(1'h0)] reg340 = (1'h0);
  reg [(3'h7):(1'h0)] reg339 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar338 = (1'h0);
  reg [(5'h11):(1'h0)] forvar337 = (1'h0);
  reg [(5'h13):(1'h0)] reg336 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg335 = (1'h0);
  reg [(3'h4):(1'h0)] reg334 = (1'h0);
  reg [(5'h13):(1'h0)] reg333 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire332;
  wire [(5'h10):(1'h0)] wire331;
  reg signed [(5'h15):(1'h0)] reg330 = (1'h0);
  reg [(5'h13):(1'h0)] reg329 = (1'h0);
  reg [(4'he):(1'h0)] reg328 = (1'h0);
  reg [(5'h15):(1'h0)] reg327 = (1'h0);
  reg [(4'h8):(1'h0)] reg326 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg325 = (1'h0);
  reg [(3'h5):(1'h0)] forvar324 = (1'h0);
  reg [(2'h3):(1'h0)] reg323 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg322 = (1'h0);
  reg [(2'h2):(1'h0)] reg321 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar320 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg319 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg318 = (1'h0);
  wire [(3'h5):(1'h0)] wire317;
  wire [(5'h10):(1'h0)] wire316;
  wire signed [(4'ha):(1'h0)] wire315;
  reg [(4'h9):(1'h0)] reg314 = (1'h0);
  reg [(3'h6):(1'h0)] reg313 = (1'h0);
  reg [(4'he):(1'h0)] reg312 = (1'h0);
  reg [(5'h12):(1'h0)] reg311 = (1'h0);
  reg [(5'h12):(1'h0)] reg310 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar309 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg308 = (1'h0);
  wire [(4'h9):(1'h0)] wire307;
  wire [(5'h14):(1'h0)] wire306;
  wire [(4'hb):(1'h0)] wire305;
  wire [(3'h4):(1'h0)] wire304;
  reg [(2'h2):(1'h0)] reg303 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg302 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg301 = (1'h0);
  reg [(3'h5):(1'h0)] reg300 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg299 = (1'h0);
  reg [(4'he):(1'h0)] reg298 = (1'h0);
  reg [(5'h10):(1'h0)] reg297 = (1'h0);
  reg [(4'hc):(1'h0)] reg296 = (1'h0);
  reg [(5'h14):(1'h0)] forvar295 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg294 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg293 = (1'h0);
  reg [(4'hf):(1'h0)] forvar292 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg291 = (1'h0);
  wire [(3'h5):(1'h0)] wire290;
  assign y = {wire347,
                 wire346,
                 reg345,
                 reg344,
                 reg343,
                 reg342,
                 reg341,
                 reg340,
                 reg339,
                 forvar338,
                 forvar337,
                 reg336,
                 reg335,
                 reg334,
                 reg333,
                 wire332,
                 wire331,
                 reg330,
                 reg329,
                 reg328,
                 reg327,
                 reg326,
                 reg325,
                 forvar324,
                 reg323,
                 reg322,
                 reg321,
                 forvar320,
                 reg319,
                 reg318,
                 wire317,
                 wire316,
                 wire315,
                 reg314,
                 reg313,
                 reg312,
                 reg311,
                 reg310,
                 forvar309,
                 reg308,
                 wire307,
                 wire306,
                 wire305,
                 wire304,
                 reg303,
                 reg302,
                 reg301,
                 reg300,
                 reg299,
                 reg298,
                 reg297,
                 reg296,
                 forvar295,
                 reg294,
                 reg293,
                 forvar292,
                 reg291,
                 wire290,
                 (1'h0)};
  assign wire290 = wire288;
  always
    @(posedge clk) begin
      reg291 <= wire287[(4'hc):(1'h0)];
    end
  always
    @(posedge clk) begin
      for (forvar292 = (1'h0); (forvar292 < (1'h1)); forvar292 = (forvar292 + (1'h1)))
        begin
          reg293 <= $unsigned((wire290[(3'h5):(3'h5)] ?
              (wire289 ?
                  (wire288 ?
                      (wire286 ?
                          wire286 : wire290) : wire290) : $unsigned((wire290 ?
                      wire290 : (8'hb1)))) : forvar292));
          reg294 <= (reg291 ?
              (((8'hbb) ?
                  wire290[(2'h2):(2'h2)] : reg293[(5'h11):(3'h7)]) * ((~((8'ha8) ?
                  wire286 : forvar292)) && (((8'hb3) | wire286) && wire288))) : wire290[(3'h4):(2'h3)]);
          for (forvar295 = (1'h0); (forvar295 < (1'h1)); forvar295 = (forvar295 + (1'h1)))
            begin
              reg296 <= wire287[(4'hd):(4'ha)];
              reg297 <= (wire286[(1'h0):(1'h0)] <<< reg293[(4'hd):(4'hd)]);
              reg298 = (|$unsigned($unsigned({$unsigned(wire287),
                  (|wire290)})));
            end
          reg299 <= (^~reg293[(4'hb):(3'h5)]);
        end
      reg300 <= $unsigned(reg298[(3'h7):(1'h1)]);
      reg301 <= wire288[(3'h6):(3'h6)];
      reg302 <= {$unsigned(reg296[(3'h5):(2'h3)])};
      reg303 <= $unsigned(reg301[(4'hf):(4'h8)]);
    end
  assign wire304 = wire288[(2'h2):(2'h2)];
  assign wire305 = reg293;
  assign wire306 = (&{{$unsigned((|reg293))}});
  assign wire307 = (wire288 <= reg297);
  always
    @(posedge clk) begin
      reg308 <= ((wire304[(3'h4):(2'h3)] ^ ($unsigned($unsigned(reg303)) ?
              (^~(reg291 >>> reg300)) : (reg293[(2'h2):(2'h2)] * (^~(8'ha8))))) ?
          reg303 : wire305[(3'h4):(2'h2)]);
      for (forvar309 = (1'h0); (forvar309 < (2'h3)); forvar309 = (forvar309 + (1'h1)))
        begin
          reg310 = forvar295;
          reg311 <= ((reg310 != (-(wire304[(1'h0):(1'h0)] <<< $signed(forvar295)))) ?
              {($signed((reg310 ?
                      forvar309 : wire307)) >>> wire286)} : {reg293});
        end
      reg312 <= (((((+wire288) <= reg294[(3'h6):(3'h5)]) ?
          $signed((reg297 ?
              wire287 : (8'ha9))) : ($unsigned(reg297) * reg294[(3'h6):(3'h4)])) - $signed(reg293[(4'hc):(2'h3)])) ^ $signed(((8'hb5) >= $unsigned(wire304))));
      reg313 <= ((^~reg294[(3'h7):(2'h2)]) == ($signed(reg297[(3'h7):(2'h2)]) >> $unsigned($signed((~|(8'hb1))))));
      reg314 <= {(7'h40)};
    end
  assign wire315 = $signed((wire290 >> $unsigned(wire306)));
  assign wire316 = ($signed((wire307 == reg296[(1'h0):(1'h0)])) ^ $unsigned((8'ha8)));
  assign wire317 = {{$signed($unsigned($unsigned(wire286)))},
                       ((reg312[(1'h0):(1'h0)] ? reg302 : $signed(reg296)) ?
                           $signed(wire289) : {(reg311[(4'h8):(4'h8)] ?
                                   reg296 : forvar292[(3'h4):(2'h2)])})};
  always
    @(posedge clk) begin
      reg318 = $unsigned($unsigned($unsigned((~|(^~wire306)))));
      reg319 <= (+(~|$unsigned($signed(reg308[(3'h6):(3'h5)]))));
    end
  always
    @(posedge clk) begin
      for (forvar320 = (1'h0); (forvar320 < (3'h4)); forvar320 = (forvar320 + (1'h1)))
        begin
          reg321 = ($signed($signed((reg310 >> $unsigned(reg303)))) >> reg300[(2'h2):(1'h1)]);
          reg322 <= (((forvar320[(3'h5):(2'h3)] ?
              forvar292 : reg301) << (wire287 ?
              reg291[(3'h5):(2'h2)] : $signed($unsigned(wire307)))) >= (((!(~^reg314)) && (^$unsigned(reg302))) - wire316));
        end
      reg323 <= {(7'h40), $signed((^$signed({wire316})))};
      for (forvar324 = (1'h0); (forvar324 < (1'h1)); forvar324 = (forvar324 + (1'h1)))
        begin
          reg325 <= reg308[(3'h6):(3'h4)];
          reg326 <= $unsigned((reg310[(3'h7):(2'h3)] ?
              $signed(reg297[(1'h0):(1'h0)]) : $unsigned(reg308[(3'h4):(1'h1)])));
          reg327 <= wire304;
          reg328 = reg311;
          reg329 = (^~(!reg300[(1'h0):(1'h0)]));
        end
    end
  always
    @(posedge clk) begin
      reg330 <= $signed(wire315);
    end
  assign wire331 = $unsigned(reg310[(4'h9):(2'h2)]);
  assign wire332 = forvar295[(5'h11):(4'hd)];
  always
    @(posedge clk) begin
      reg333 <= {($unsigned($unsigned($signed((8'hb7)))) - $unsigned(wire332[(4'h8):(2'h2)]))};
      reg334 <= (((^~(((8'hbb) - (8'ha5)) ?
                  (wire305 ? wire304 : reg303) : $unsigned(reg298))) ?
              $signed($unsigned((reg293 ? reg325 : reg325))) : reg330) ?
          reg326 : ({$signed((reg329 ? forvar295 : reg302)), reg313} ?
              (~^((reg293 == (8'hb1)) ?
                  $unsigned(wire316) : $signed(forvar324))) : $unsigned(reg296)));
      reg335 <= {({reg321[(1'h0):(1'h0)]} ?
              {$unsigned(reg321)} : $signed(($unsigned(wire315) < wire331)))};
      reg336 = $unsigned($signed($unsigned($signed($unsigned(reg296)))));
      for (forvar337 = (1'h0); (forvar337 < (2'h2)); forvar337 = (forvar337 + (1'h1)))
        begin
          for (forvar338 = (1'h0); (forvar338 < (2'h2)); forvar338 = (forvar338 + (1'h1)))
            begin
              reg339 <= $signed(((^(forvar324[(2'h2):(1'h0)] >= (~(8'hb0)))) ?
                  (((wire289 ? wire289 : reg302) >>> (wire332 <<< wire304)) ?
                      ($unsigned(wire288) ?
                          forvar309 : (wire288 ?
                              reg297 : (8'hb8))) : reg297) : ($signed((+reg311)) ?
                      {$signed(wire287)} : $signed(reg308[(3'h4):(2'h3)]))));
              reg340 <= (-$unsigned((!forvar337)));
              reg341 <= {(-(-(&reg296[(2'h2):(2'h2)]))),
                  (wire287[(4'h8):(4'h8)] ?
                      ($unsigned(forvar292[(4'hb):(3'h4)]) >>> forvar320[(3'h5):(1'h1)]) : {(8'hb5),
                          $signed(reg291[(2'h3):(2'h2)])})};
              reg342 <= (^$unsigned((|(reg308[(1'h1):(1'h0)] > $unsigned(reg336)))));
            end
          reg343 <= $unsigned(((8'h9f) == wire290[(2'h2):(1'h0)]));
          reg344 <= {forvar292[(4'hf):(3'h5)],
              $unsigned($signed(((~|reg334) <= (reg303 ? reg340 : reg327))))};
          reg345 <= $signed((~reg342));
        end
    end
  assign wire346 = wire304[(2'h2):(1'h1)];
  assign wire347 = $unsigned(({$unsigned(reg336[(2'h3):(1'h0)]),
                       reg334} < $signed((!(8'ha2)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module111  (y, clk, wire112, wire113, wire114, wire115);
  output wire [(32'h49):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire112;
  input wire [(5'h13):(1'h0)] wire113;
  input wire signed [(5'h13):(1'h0)] wire114;
  input wire signed [(4'hd):(1'h0)] wire115;
  reg [(3'h5):(1'h0)] reg277 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg276 = (1'h0);
  reg [(3'h5):(1'h0)] reg275 = (1'h0);
  wire [(5'h13):(1'h0)] wire274;
  wire [(5'h11):(1'h0)] wire273;
  wire signed [(4'hb):(1'h0)] wire116;
  wire [(3'h7):(1'h0)] wire271;
  assign y = {reg277,
                 reg276,
                 reg275,
                 wire274,
                 wire273,
                 wire116,
                 wire271,
                 (1'h0)};
  assign wire116 = $unsigned(wire112);
  module117 modinst272 (wire271, clk, wire115, wire114, wire112, wire116, wire113);
  assign wire273 = {$unsigned({wire115,
                           ((wire113 >>> wire116) ^~ $signed(wire116))})};
  assign wire274 = (wire271[(3'h7):(2'h2)] <= ($signed({((8'hb3) ^ (8'had)),
                       $unsigned(wire116)}) < (^~wire116[(1'h1):(1'h0)])));
  always
    @(posedge clk) begin
      reg275 <= ((wire271[(3'h4):(3'h4)] ^ ({(wire112 ?
              (8'hbf) : wire114)} ^ $unsigned({wire114}))) > wire113);
      reg276 <= ($unsigned(wire274[(3'h4):(3'h4)]) ?
          $signed(wire115[(4'h9):(3'h5)]) : $signed(($unsigned((wire115 >= (8'hb6))) ?
              ((!(8'hb8)) ^ wire116) : ((8'ha7) ?
                  ((8'hb4) ? reg275 : wire273) : ((8'ha2) >>> wire116)))));
      reg277 <= (reg276[(4'h8):(1'h1)] ?
          {{reg276[(3'h7):(3'h4)]},
              wire115} : $signed($signed($unsigned($unsigned(wire112)))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module83
#( parameter param100 = ((((((8'h9e) > (8'ha9)) ? (~^(8'haa)) : ((8'ha2) ^~ (8'ha0))) ? (8'hb7) : (+(+(8'hb5)))) ? {({(8'hb1), (8'ha2)} ? ((8'ha6) ? (8'hb9) : (8'hbc)) : (~|(8'ha5))), (7'h41)} : ((((8'hbc) < (8'haa)) == ((8'hb9) ^~ (8'h9c))) > {((7'h41) == (7'h44)), ((8'haa) >= (8'ha1))})) ? ((((~|(7'h41)) ? ((8'hb3) >>> (8'hba)) : ((8'ha7) + (8'h9c))) ? (((8'hbf) >> (7'h44)) ? ((8'hb5) ^~ (8'ha8)) : {(7'h42)}) : (((8'h9d) ? (8'h9e) : (8'hba)) ~^ ((8'ha3) ? (8'hbf) : (7'h43)))) ? {(((8'hb0) ~^ (8'h9c)) ? ((8'hac) ? (8'hbc) : (8'hac)) : ((8'hac) ? (7'h43) : (8'hae))), ({(8'hb2), (8'h9d)} != ((8'ha4) ? (8'ha2) : (8'ha9)))} : ({((8'hae) & (8'hb0)), (8'ha2)} && ((~|(8'hbc)) >>> ((8'hb3) ? (8'ha4) : (8'hb0))))) : (+(((&(7'h42)) ? ((7'h43) ^~ (8'hb5)) : ((8'haf) << (8'ha7))) ~^ (8'ha0)))) )
(y, clk, wire88, wire87, wire86, wire85, wire84);
  output wire [(32'h6c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h9):(1'h0)] wire88;
  input wire [(4'hf):(1'h0)] wire87;
  input wire signed [(3'h5):(1'h0)] wire86;
  input wire signed [(4'ha):(1'h0)] wire85;
  input wire [(4'h9):(1'h0)] wire84;
  reg [(2'h3):(1'h0)] reg99 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire98;
  reg signed [(4'hc):(1'h0)] reg97 = (1'h0);
  reg [(5'h11):(1'h0)] reg96 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg95 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg94 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar93 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg92 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg91 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire90;
  wire signed [(4'h8):(1'h0)] wire89;
  assign y = {reg99,
                 wire98,
                 reg97,
                 reg96,
                 reg95,
                 reg94,
                 forvar93,
                 reg92,
                 reg91,
                 wire90,
                 wire89,
                 (1'h0)};
  assign wire89 = wire88;
  assign wire90 = wire89;
  always
    @(posedge clk) begin
      reg91 <= $unsigned(wire89);
      reg92 <= wire84[(2'h3):(1'h1)];
      for (forvar93 = (1'h0); (forvar93 < (1'h0)); forvar93 = (forvar93 + (1'h1)))
        begin
          reg94 = (wire88[(3'h6):(3'h5)] ?
              (((reg91 < ((8'ha0) ? reg92 : (7'h41))) ?
                  $unsigned($signed(wire87)) : ((wire90 ?
                      wire88 : wire85) ~^ (-wire87))) || (({reg91,
                      wire88} <= {wire88, wire87}) ?
                  (wire85[(3'h7):(1'h0)] ?
                      wire86[(3'h4):(1'h0)] : $unsigned(forvar93)) : ((!(8'had)) ?
                      $unsigned(reg91) : wire89[(2'h2):(1'h0)]))) : $signed(forvar93));
          reg95 <= (wire84 ? (8'hb5) : wire89[(1'h0):(1'h0)]);
        end
      reg96 = reg95[(2'h2):(1'h0)];
      reg97 = (forvar93 < (|$signed($signed((~^reg92)))));
    end
  assign wire98 = ((~&{((~^reg92) ? reg97 : $unsigned(forvar93)),
                          ((^~wire89) + (|wire90))}) ?
                      $unsigned(({((8'h9e) >>> reg91)} ?
                          $signed($unsigned(reg97)) : (|(|wire90)))) : wire86);
  always
    @(posedge clk) begin
      reg99 <= wire85[(1'h0):(1'h0)];
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module117
#( parameter param270 = ((^~((((8'ha1) ? (8'haa) : (8'h9f)) && ((8'hb1) >>> (8'ha2))) <= (~&(~^(8'hab))))) ? (!((((8'hac) ? (7'h42) : (8'hb3)) + (!(8'had))) ? {(8'ha5), (&(8'hac))} : (~(|(8'hbe))))) : (~^{(8'ha5)})) )
(y, clk, wire122, wire121, wire120, wire119, wire118);
  output wire [(32'hf3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h7):(1'h0)] wire122;
  input wire signed [(2'h2):(1'h0)] wire121;
  input wire [(5'h14):(1'h0)] wire120;
  input wire signed [(3'h5):(1'h0)] wire119;
  input wire [(5'h13):(1'h0)] wire118;
  wire [(5'h11):(1'h0)] wire183;
  reg [(4'he):(1'h0)] reg137 = (1'h0);
  reg [(4'hc):(1'h0)] reg136 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg135 = (1'h0);
  wire [(4'hc):(1'h0)] wire134;
  reg [(4'hf):(1'h0)] reg133 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg132 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg131 = (1'h0);
  wire [(5'h11):(1'h0)] wire130;
  reg signed [(4'hd):(1'h0)] reg129 = (1'h0);
  reg [(4'hd):(1'h0)] reg128 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg127 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg126 = (1'h0);
  wire [(5'h12):(1'h0)] wire125;
  wire [(5'h13):(1'h0)] wire124;
  reg [(2'h2):(1'h0)] reg123 = (1'h0);
  wire [(4'hc):(1'h0)] wire185;
  wire [(3'h7):(1'h0)] wire268;
  assign y = {wire183,
                 reg137,
                 reg136,
                 reg135,
                 wire134,
                 reg133,
                 reg132,
                 reg131,
                 wire130,
                 reg129,
                 reg128,
                 reg127,
                 reg126,
                 wire125,
                 wire124,
                 reg123,
                 wire185,
                 wire268,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg123 <= (((wire119 ? (~^$signed(wire119)) : (wire121 | wire120)) ?
          wire119 : (wire121 ^~ $signed($unsigned(wire120)))) != $unsigned(wire121));
    end
  assign wire124 = wire119[(3'h4):(2'h2)];
  assign wire125 = $signed(((~^$unsigned((!wire118))) ?
                       $signed($unsigned(wire120[(4'h9):(4'h8)])) : wire119));
  always
    @(posedge clk) begin
      reg126 <= {$signed($signed(({wire121} ? wire124 : (^~(8'hb6))))),
          wire122};
      reg127 <= $unsigned(((~|($signed(wire125) + {wire119})) ^ (^wire118[(4'hd):(4'h9)])));
      reg128 <= (((wire119 ?
              $signed((reg123 ? wire122 : reg127)) : (((8'ha8) ?
                  wire122 : wire121) - $unsigned(reg126))) ?
          ($unsigned($signed(reg123)) ?
              wire124 : wire121) : wire125) - $signed(($unsigned((wire121 ?
          reg127 : wire121)) <= wire119)));
      reg129 <= ($unsigned({(!$unsigned((7'h43))), wire124[(4'ha):(4'h9)]}) ?
          $signed(((wire122[(3'h7):(2'h3)] ?
                  $signed(wire118) : $unsigned(wire119)) ?
              {$signed(wire125)} : wire120[(4'hb):(4'h9)])) : ($signed(((wire119 || wire118) < (wire124 ?
              wire120 : wire121))) <= (~$unsigned((|reg123)))));
    end
  assign wire130 = $unsigned($unsigned({(!((7'h42) ^~ wire119)),
                       {$signed(wire119), (reg129 | wire120)}}));
  always
    @(posedge clk) begin
      reg131 = wire124[(2'h2):(2'h2)];
      reg132 = (((wire130 >> (wire125 || {wire130})) << reg129) << $signed({(~|reg123[(1'h1):(1'h0)])}));
      reg133 <= $unsigned($signed(($unsigned($unsigned((7'h41))) ?
          ($unsigned(reg127) ?
              {wire125} : ((8'haa) - reg128)) : $unsigned((wire121 ?
              wire124 : reg123)))));
    end
  assign wire134 = {wire122[(2'h2):(1'h0)],
                       ((wire121 ?
                           (8'hb4) : {$unsigned(wire119)}) <= $signed(($signed(reg123) && (wire118 ?
                           reg128 : wire118))))};
  always
    @(posedge clk) begin
      reg135 <= $unsigned(wire121[(2'h2):(2'h2)]);
      reg136 <= $signed(wire121[(1'h0):(1'h0)]);
      reg137 <= wire130[(4'h9):(3'h6)];
    end
  module138 modinst184 (.clk(clk), .wire139(reg126), .y(wire183), .wire141(reg129), .wire143(reg132), .wire142(reg137), .wire140(wire124));
  assign wire185 = $signed($unsigned((^~((reg129 ?
                       reg135 : wire122) & $unsigned(wire119)))));
  module186 modinst269 (.clk(clk), .wire188(wire120), .wire191(wire134), .wire189(reg133), .wire187(reg131), .wire190(reg135), .y(wire268));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module186
#(parameter param267 = (~(^~(&(~|((8'hb6) ? (8'hbe) : (8'hbd)))))))
(y, clk, wire191, wire190, wire189, wire188, wire187);
  output wire [(32'h36d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire191;
  input wire [(5'h11):(1'h0)] wire190;
  input wire [(4'hf):(1'h0)] wire189;
  input wire signed [(5'h14):(1'h0)] wire188;
  input wire [(5'h15):(1'h0)] wire187;
  reg signed [(4'hd):(1'h0)] reg266 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg265 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg264 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire263;
  reg [(5'h11):(1'h0)] reg262 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg261 = (1'h0);
  reg [(3'h7):(1'h0)] reg260 = (1'h0);
  reg [(4'h9):(1'h0)] reg259 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg258 = (1'h0);
  reg [(5'h14):(1'h0)] reg257 = (1'h0);
  reg [(5'h10):(1'h0)] forvar256 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg255 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg254 = (1'h0);
  reg [(5'h14):(1'h0)] reg253 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg252 = (1'h0);
  reg [(4'hc):(1'h0)] reg251 = (1'h0);
  reg [(3'h6):(1'h0)] reg250 = (1'h0);
  reg [(4'h9):(1'h0)] reg249 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg248 = (1'h0);
  reg [(5'h14):(1'h0)] reg247 = (1'h0);
  reg [(4'he):(1'h0)] reg246 = (1'h0);
  reg [(4'ha):(1'h0)] reg245 = (1'h0);
  reg signed [(4'he):(1'h0)] reg244 = (1'h0);
  reg [(3'h6):(1'h0)] reg243 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg242 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar241 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg240 = (1'h0);
  reg [(4'h9):(1'h0)] forvar239 = (1'h0);
  reg [(4'ha):(1'h0)] reg238 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg237 = (1'h0);
  reg [(2'h2):(1'h0)] reg236 = (1'h0);
  reg [(5'h11):(1'h0)] reg235 = (1'h0);
  reg [(4'hd):(1'h0)] reg234 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg233 = (1'h0);
  reg [(3'h4):(1'h0)] reg232 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire231;
  reg signed [(3'h7):(1'h0)] reg230 = (1'h0);
  reg [(4'he):(1'h0)] reg229 = (1'h0);
  reg [(4'h8):(1'h0)] reg228 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg227 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg226 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg225 = (1'h0);
  wire [(3'h6):(1'h0)] wire224;
  wire signed [(4'hc):(1'h0)] wire223;
  reg [(5'h10):(1'h0)] reg222 = (1'h0);
  reg [(2'h3):(1'h0)] reg221 = (1'h0);
  reg [(4'he):(1'h0)] reg220 = (1'h0);
  reg [(5'h10):(1'h0)] reg219 = (1'h0);
  reg [(5'h12):(1'h0)] reg218 = (1'h0);
  reg [(3'h4):(1'h0)] reg217 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg216 = (1'h0);
  reg [(4'h8):(1'h0)] forvar215 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg214 = (1'h0);
  reg [(3'h5):(1'h0)] reg213 = (1'h0);
  reg [(3'h4):(1'h0)] reg212 = (1'h0);
  reg [(5'h15):(1'h0)] reg211 = (1'h0);
  reg [(3'h6):(1'h0)] forvar210 = (1'h0);
  reg [(5'h11):(1'h0)] reg210 = (1'h0);
  reg [(3'h5):(1'h0)] reg209 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg208 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg207 = (1'h0);
  reg [(4'he):(1'h0)] reg206 = (1'h0);
  reg [(3'h7):(1'h0)] reg205 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg204 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg203 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar202 = (1'h0);
  reg signed [(4'he):(1'h0)] reg201 = (1'h0);
  reg [(4'he):(1'h0)] reg200 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg199 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar198 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg197 = (1'h0);
  reg [(4'hf):(1'h0)] forvar196 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg195 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg194 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg193 = (1'h0);
  reg [(5'h13):(1'h0)] reg192 = (1'h0);
  assign y = {reg266,
                 reg265,
                 reg264,
                 wire263,
                 reg262,
                 reg261,
                 reg260,
                 reg259,
                 reg258,
                 reg257,
                 forvar256,
                 reg255,
                 reg254,
                 reg253,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 reg248,
                 reg247,
                 reg246,
                 reg245,
                 reg244,
                 reg243,
                 reg242,
                 forvar241,
                 reg240,
                 forvar239,
                 reg238,
                 reg237,
                 reg236,
                 reg235,
                 reg234,
                 reg233,
                 reg232,
                 wire231,
                 reg230,
                 reg229,
                 reg228,
                 reg227,
                 reg226,
                 reg225,
                 wire224,
                 wire223,
                 reg222,
                 reg221,
                 reg220,
                 reg219,
                 reg218,
                 reg217,
                 reg216,
                 forvar215,
                 reg214,
                 reg213,
                 reg212,
                 reg211,
                 forvar210,
                 reg210,
                 reg209,
                 reg208,
                 reg207,
                 reg206,
                 reg205,
                 reg204,
                 reg203,
                 forvar202,
                 reg201,
                 reg200,
                 reg199,
                 forvar198,
                 reg197,
                 forvar196,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg192 <= wire187;
      reg193 = ({(|{(wire191 ? wire189 : reg192)})} ?
          (~&(|wire189[(4'hc):(4'hc)])) : $signed(reg192[(3'h7):(2'h2)]));
      reg194 <= ($signed(((8'hb4) ?
          reg193[(3'h4):(1'h0)] : wire187)) | (reg192 | ({{(7'h42)}} ?
          ((wire189 * (8'haf)) + (wire191 ?
              (8'hb3) : wire190)) : (!$unsigned(wire189)))));
      reg195 = $unsigned($signed(wire189[(4'hc):(3'h7)]));
    end
  always
    @(posedge clk) begin
      for (forvar196 = (1'h0); (forvar196 < (2'h3)); forvar196 = (forvar196 + (1'h1)))
        begin
          reg197 <= ((8'hbb) ?
              ((8'hb0) | ($signed(wire190) ?
                  reg195[(1'h0):(1'h0)] : $signed($unsigned((7'h44))))) : $signed((^~{wire187})));
          for (forvar198 = (1'h0); (forvar198 < (1'h0)); forvar198 = (forvar198 + (1'h1)))
            begin
              reg199 <= reg195[(3'h6):(3'h5)];
              reg200 <= ((({$signed(reg199),
                      $signed(reg197)} - $signed((wire187 < wire191))) <= reg197) ?
                  ($signed(wire187) ?
                      {(!$signed((8'hb9)))} : $unsigned(((reg193 >> reg197) ?
                          {reg194,
                              wire189} : $unsigned(reg195)))) : $unsigned((|{reg197,
                      $signed(wire189)})));
            end
          reg201 <= (8'hb1);
          for (forvar202 = (1'h0); (forvar202 < (1'h0)); forvar202 = (forvar202 + (1'h1)))
            begin
              reg203 = ((&reg200[(1'h1):(1'h1)]) + $unsigned((~&((|wire191) ?
                  wire187[(3'h4):(2'h3)] : $signed(reg199)))));
              reg204 <= ($signed(reg201) >> {(~&(~|(reg195 ^~ wire187))),
                  $signed(((wire189 || wire188) ?
                      {reg193, wire189} : (reg192 >> reg193)))});
              reg205 = wire188;
              reg206 <= {$signed(wire187[(5'h15):(1'h0)])};
              reg207 = forvar202[(5'h11):(4'hb)];
            end
          reg208 <= (~|$signed((8'haa)));
        end
      if ((^~$unsigned(reg199)))
        begin
          reg209 = {{$unsigned((~^(reg197 == wire187)))}};
          reg210 <= (&($unsigned($unsigned($unsigned(reg208))) ?
              forvar198[(2'h3):(2'h3)] : {(wire187[(4'hc):(4'h8)] ^ reg204[(3'h5):(2'h3)]),
                  $signed($unsigned(reg200))}));
        end
      else
        begin
          reg209 <= (-reg194);
          for (forvar210 = (1'h0); (forvar210 < (2'h3)); forvar210 = (forvar210 + (1'h1)))
            begin
              reg211 <= {$signed(forvar210)};
              reg212 <= $signed($unsigned((8'hb3)));
              reg213 <= $unsigned(reg195[(1'h0):(1'h0)]);
              reg214 = (&reg195[(1'h0):(1'h0)]);
            end
          for (forvar215 = (1'h0); (forvar215 < (1'h0)); forvar215 = (forvar215 + (1'h1)))
            begin
              reg216 <= reg209[(3'h5):(2'h2)];
              reg217 = reg212[(2'h3):(2'h2)];
              reg218 = (~((!forvar215) <<< ((8'ha1) & forvar210[(3'h5):(2'h2)])));
              reg219 <= ($unsigned(((+(-forvar198)) ?
                  (|((8'hbb) <<< reg218)) : ((forvar196 ? reg201 : forvar210) ?
                      reg199 : (reg212 ?
                          reg193 : reg201)))) <<< (~^$signed(($unsigned(forvar210) ^ (reg197 | reg193)))));
            end
        end
      reg220 <= reg217;
      reg221 <= ($unsigned(reg208[(3'h4):(2'h2)]) & $signed($unsigned(reg219[(4'he):(3'h7)])));
      reg222 <= $signed(({reg204} >> reg203[(4'hb):(3'h4)]));
    end
  assign wire223 = ((^~$signed($signed({reg201}))) ~^ $unsigned(((reg197[(1'h0):(1'h0)] ?
                           reg218[(1'h1):(1'h1)] : reg206) ?
                       $unsigned($unsigned(reg212)) : ((reg197 >= reg195) > (reg222 | reg200)))));
  assign wire224 = (^~(~(reg220 | $unsigned((~^(8'hbb))))));
  always
    @(posedge clk) begin
      reg225 <= $signed((forvar198[(2'h3):(1'h1)] ?
          $unsigned(reg192) : $unsigned(wire187[(5'h13):(3'h4)])));
    end
  always
    @(posedge clk) begin
      reg226 <= ($signed($unsigned(($signed(reg220) >>> $signed((8'hbe))))) << $unsigned((reg210 ?
          reg201 : $signed($unsigned(reg193)))));
      reg227 <= ({$signed($signed((-reg208))),
          $unsigned({$signed(reg226), (8'hb6)})} ^~ ({(7'h42),
              (^(reg226 ? reg220 : (8'hb9)))} ?
          (wire190 ?
              $unsigned($unsigned(wire190)) : ((forvar196 & reg204) != (-(8'hab)))) : $unsigned($unsigned((reg214 ?
              reg201 : reg214)))));
      reg228 <= ((~^(reg210 * (wire191 <<< (wire189 ? reg205 : reg199)))) ?
          (~^$signed((~&reg213))) : ($unsigned(reg216) ?
              $unsigned({$unsigned((8'hbe)), (~^reg210)}) : reg194));
      reg229 <= (|$signed(reg221));
      reg230 <= (8'hba);
    end
  assign wire231 = ($unsigned(wire190) ?
                       (8'hac) : $signed(((8'hb7) ?
                           ((reg203 != reg218) >= (reg214 ?
                               forvar198 : reg199)) : forvar210[(1'h1):(1'h0)])));
  always
    @(posedge clk) begin
      reg232 <= $unsigned((!({(reg217 || reg199)} == $signed($signed(reg225)))));
      reg233 = forvar215;
      reg234 <= reg205;
      reg235 <= $signed((~^wire189));
    end
  always
    @(posedge clk) begin
      reg236 <= (((8'h9f) ?
              $unsigned((~{(7'h43), (8'hb3)})) : ($signed($signed((8'hb7))) ?
                  $unsigned({reg211}) : ((wire224 ? reg230 : reg216) ?
                      wire223 : (reg227 * reg225)))) ?
          reg230 : $signed((forvar202 ?
              (~|$unsigned(reg203)) : $unsigned($signed(wire224)))));
      reg237 <= $signed(reg194);
      reg238 <= (^forvar215);
      for (forvar239 = (1'h0); (forvar239 < (1'h0)); forvar239 = (forvar239 + (1'h1)))
        begin
          reg240 <= (~$signed($unsigned($unsigned({wire231, reg216}))));
          for (forvar241 = (1'h0); (forvar241 < (2'h3)); forvar241 = (forvar241 + (1'h1)))
            begin
              reg242 <= ($unsigned((($signed(reg229) ?
                          $unsigned(forvar239) : {reg193}) ?
                      wire231 : reg220[(4'h9):(3'h7)])) ?
                  ((8'hbd) ?
                      reg228[(3'h6):(2'h3)] : reg237) : (~(($unsigned(reg210) ?
                          ((8'hbc) || reg214) : $signed(reg229)) ?
                      (forvar202[(1'h0):(1'h0)] ?
                          $signed(reg225) : $unsigned(reg227)) : $unsigned(reg222[(3'h4):(1'h1)]))));
              reg243 = reg237[(5'h12):(3'h6)];
              reg244 <= $signed(reg234[(4'h9):(3'h4)]);
              reg245 = $unsigned({reg236});
              reg246 = (reg194[(4'hb):(2'h2)] & $unsigned(reg225));
            end
          reg247 <= $signed($unsigned(reg222[(4'he):(4'hb)]));
        end
    end
  always
    @(posedge clk) begin
      reg248 <= (-reg226[(1'h0):(1'h0)]);
      reg249 <= reg204;
      reg250 <= reg207;
    end
  always
    @(posedge clk) begin
      reg251 <= $unsigned(wire231[(2'h3):(2'h3)]);
      reg252 <= wire188;
      reg253 = (reg207[(3'h5):(2'h3)] & {reg238[(2'h3):(2'h2)],
          $unsigned($unsigned((reg209 * reg220)))});
      reg254 <= (($unsigned((reg201[(2'h2):(2'h2)] ?
              (reg235 >>> (8'ha5)) : (reg217 || reg230))) ?
          (^~$unsigned(wire189[(2'h2):(1'h0)])) : (-{((8'ha8) >> reg246),
              reg250})) ^ reg192[(4'h8):(2'h3)]);
    end
  always
    @(posedge clk) begin
      reg255 = wire187;
      for (forvar256 = (1'h0); (forvar256 < (1'h0)); forvar256 = (forvar256 + (1'h1)))
        begin
          reg257 <= reg234;
          reg258 = $signed($unsigned($signed((8'hb6))));
          reg259 <= (&reg213[(2'h3):(2'h3)]);
        end
      reg260 = reg213[(1'h0):(1'h0)];
      reg261 <= ((((forvar215 ?
              reg203 : (^~wire224)) <= ({reg246} && $signed(reg225))) >>> {((reg221 | reg237) != (reg257 ?
                  (8'hb2) : reg250)),
              $unsigned(reg209[(1'h0):(1'h0)])}) ?
          $unsigned(reg244[(1'h0):(1'h0)]) : $signed(reg259[(1'h0):(1'h0)]));
      reg262 <= (8'ha1);
    end
  assign wire263 = (~(8'ha6));
  always
    @(posedge clk) begin
      reg264 = ((~&$signed((((8'had) ? forvar256 : (8'ha4)) && ((8'h9e) ?
              reg201 : (8'hb6))))) ?
          (&(|$signed((!(8'hb3))))) : reg247);
      reg265 <= reg216[(2'h2):(2'h2)];
      reg266 = reg253[(4'h8):(2'h3)];
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module138  (y, clk, wire143, wire142, wire141, wire140, wire139);
  output wire [(32'h1b4):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire143;
  input wire [(4'h9):(1'h0)] wire142;
  input wire signed [(4'h9):(1'h0)] wire141;
  input wire signed [(5'h13):(1'h0)] wire140;
  input wire [(4'hb):(1'h0)] wire139;
  reg [(5'h15):(1'h0)] reg182 = (1'h0);
  reg [(4'h8):(1'h0)] reg181 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg180 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg179 = (1'h0);
  reg [(4'hd):(1'h0)] reg178 = (1'h0);
  reg [(5'h15):(1'h0)] reg177 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg176 = (1'h0);
  reg [(5'h12):(1'h0)] reg175 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg174 = (1'h0);
  reg [(4'he):(1'h0)] forvar173 = (1'h0);
  reg [(5'h11):(1'h0)] reg172 = (1'h0);
  reg [(5'h10):(1'h0)] reg171 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg170 = (1'h0);
  reg [(3'h6):(1'h0)] reg169 = (1'h0);
  reg [(2'h3):(1'h0)] reg168 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar167 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar166 = (1'h0);
  reg [(4'hf):(1'h0)] reg165 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg164 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg163 = (1'h0);
  reg [(5'h13):(1'h0)] reg162 = (1'h0);
  reg [(3'h5):(1'h0)] forvar161 = (1'h0);
  reg [(4'h8):(1'h0)] reg160 = (1'h0);
  reg [(4'h9):(1'h0)] reg159 = (1'h0);
  reg [(4'h9):(1'h0)] reg158 = (1'h0);
  reg [(4'h8):(1'h0)] reg157 = (1'h0);
  reg [(5'h13):(1'h0)] reg156 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar155 = (1'h0);
  wire [(4'hb):(1'h0)] wire154;
  wire [(4'ha):(1'h0)] wire153;
  wire [(4'he):(1'h0)] wire152;
  reg signed [(3'h6):(1'h0)] reg151 = (1'h0);
  wire signed [(4'he):(1'h0)] wire150;
  reg [(4'h8):(1'h0)] reg149 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg148 = (1'h0);
  reg [(3'h6):(1'h0)] reg147 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg146 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg145 = (1'h0);
  reg [(4'he):(1'h0)] reg144 = (1'h0);
  assign y = {reg182,
                 reg181,
                 reg180,
                 reg179,
                 reg178,
                 reg177,
                 reg176,
                 reg175,
                 reg174,
                 forvar173,
                 reg172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 forvar167,
                 forvar166,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 forvar161,
                 reg160,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 forvar155,
                 wire154,
                 wire153,
                 wire152,
                 reg151,
                 wire150,
                 reg149,
                 reg148,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg144 <= $signed(wire140[(5'h12):(4'h9)]);
      reg145 = wire140;
      reg146 <= (-(wire141 ?
          (~reg145[(3'h7):(2'h2)]) : ($signed($signed(wire142)) + reg145)));
      reg147 <= (|($unsigned((~|(wire141 ?
          (8'hbc) : reg145))) >> $unsigned($signed($signed(reg146)))));
      reg148 = reg147[(2'h2):(1'h1)];
    end
  always
    @(posedge clk) begin
      reg149 = (+($unsigned(wire141) ?
          wire141 : ($signed((reg147 ?
              wire140 : reg144)) || $signed($signed(wire140)))));
    end
  assign wire150 = (~|$unsigned(reg148));
  always
    @(posedge clk) begin
      reg151 <= wire139[(3'h6):(3'h4)];
    end
  assign wire152 = (reg149 ?
                       ($unsigned(reg144) ?
                           reg144 : wire143[(1'h1):(1'h0)]) : ($unsigned((!(&wire140))) <<< ({reg149,
                           reg144} ^ $unsigned(((8'hb9) ? reg145 : reg149)))));
  assign wire153 = $signed({reg148[(4'h8):(3'h5)], reg145});
  assign wire154 = (|$unsigned((~^$signed((~reg146)))));
  always
    @(posedge clk) begin
      for (forvar155 = (1'h0); (forvar155 < (3'h4)); forvar155 = (forvar155 + (1'h1)))
        begin
          reg156 = reg148[(4'h9):(2'h3)];
          reg157 = (wire140[(4'he):(4'h9)] || (^forvar155[(4'ha):(3'h4)]));
          reg158 <= wire142;
        end
      reg159 <= (wire154 ?
          wire154[(3'h7):(3'h5)] : $unsigned(($unsigned((reg157 >>> wire139)) == $signed(wire143))));
      reg160 <= (($signed(((reg159 ~^ reg145) ?
              $signed(reg158) : (wire153 ~^ wire153))) - $signed((~&$unsigned(reg159)))) ?
          reg144 : reg151[(3'h5):(3'h4)]);
      for (forvar161 = (1'h0); (forvar161 < (2'h3)); forvar161 = (forvar161 + (1'h1)))
        begin
          reg162 <= (-({reg149} ?
              $unsigned((reg160[(3'h6):(3'h4)] >>> $unsigned(wire143))) : reg151[(1'h0):(1'h0)]));
          reg163 <= $unsigned(($signed($signed($signed(reg157))) ?
              (~&reg156) : ($unsigned((~&reg156)) + (^{(8'hb4)}))));
          reg164 <= reg162;
          reg165 <= reg157[(2'h3):(1'h1)];
        end
      for (forvar166 = (1'h0); (forvar166 < (1'h0)); forvar166 = (forvar166 + (1'h1)))
        begin
          for (forvar167 = (1'h0); (forvar167 < (2'h3)); forvar167 = (forvar167 + (1'h1)))
            begin
              reg168 <= forvar161[(1'h0):(1'h0)];
              reg169 = (((|forvar167) ?
                      (wire154 <= ((&reg160) ?
                          reg168[(2'h3):(1'h0)] : (&(8'ha0)))) : ((~|$unsigned(wire141)) ?
                          wire143[(1'h1):(1'h1)] : (((8'hbd) != reg151) ?
                              (^reg163) : (&reg159)))) ?
                  (~&{{$unsigned(forvar155), reg151[(3'h5):(3'h5)]},
                      ($unsigned(reg148) ?
                          (8'hac) : $signed(reg164))}) : reg165[(4'h9):(4'h9)]);
              reg170 = {$signed(reg146), $signed((&reg156))};
            end
        end
    end
  always
    @(posedge clk) begin
      reg171 <= ($unsigned($unsigned($unsigned($unsigned(reg163)))) ?
          wire154[(4'hb):(3'h7)] : $unsigned(((-(^wire139)) ?
              {((8'hb0) << reg169),
                  (reg165 ?
                      reg147 : reg156)} : $signed(wire140[(5'h11):(3'h4)]))));
      reg172 = (~&(~|$unsigned($signed((~&reg144)))));
      for (forvar173 = (1'h0); (forvar173 < (3'h4)); forvar173 = (forvar173 + (1'h1)))
        begin
          reg174 <= $signed(($signed(((reg170 * (8'hb7)) != (reg144 ^~ reg169))) ?
              (~($signed(forvar167) ?
                  (reg151 ?
                      reg172 : reg145) : reg146)) : {((forvar173 == forvar166) & (~|reg163)),
                  (reg149[(2'h2):(1'h1)] ? (+reg160) : (wire153 >= (7'h44)))}));
          reg175 <= reg163[(5'h10):(3'h5)];
          reg176 = reg163;
          reg177 <= $unsigned({$unsigned(($unsigned(forvar161) ?
                  $unsigned((8'haf)) : (reg169 >>> (7'h41))))});
          reg178 = (8'haf);
        end
    end
  always
    @(posedge clk) begin
      reg179 = ($unsigned(({(wire143 * (8'hbe)), reg158} ^~ (~|(forvar173 ?
              wire152 : reg157)))) ?
          $signed(((-$unsigned(reg168)) || wire140)) : (~(((^reg163) ?
                  reg147[(3'h5):(2'h3)] : (!reg176)) ?
              ($signed(reg151) || $signed((8'hbb))) : reg163[(1'h0):(1'h0)])));
      reg180 = wire143[(3'h5):(1'h0)];
      reg181 <= (~(~&$signed(($unsigned(reg177) != (forvar166 ~^ (8'haf))))));
      reg182 <= ((~^(~&$unsigned((|reg180)))) != $signed($signed(((^wire153) - (reg176 <= reg176)))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module377
#( parameter param537 = ((!((((8'hb8) >= (8'had)) ? ((8'hbd) | (8'hb5)) : (&(7'h44))) ? {{(7'h42)}} : (((8'hb3) >>> (8'hba)) * ((8'ha4) < (8'hbc))))) ? (((((8'hb1) ? (8'hb9) : (8'ha9)) ? (~&(8'hb9)) : ((8'hb5) ? (8'haa) : (8'hb5))) ? (!(|(8'hb4))) : {((8'ha7) ^~ (8'ha3)), (!(7'h42))}) | (7'h44)) : (((((7'h40) ? (8'hbf) : (8'hbd)) ? (8'hba) : ((8'hbb) ^~ (8'hb3))) > (((8'ha8) ? (7'h41) : (8'hbb)) <<< {(8'ha0)})) ? {(&((8'ha0) | (8'hb1)))} : ((|((8'hbd) <= (8'ha5))) | (!{(8'hbe)}))))
, parameter param538 = (8'haf) )
(y, clk, wire378, wire379, wire380, wire381);
  output wire [(32'h1bd):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h15):(1'h0)] wire378;
  input wire [(3'h6):(1'h0)] wire379;
  input wire [(3'h6):(1'h0)] wire380;
  input wire signed [(4'hc):(1'h0)] wire381;
  wire signed [(3'h5):(1'h0)] wire535;
  wire [(5'h15):(1'h0)] wire455;
  wire signed [(4'ha):(1'h0)] wire454;
  wire signed [(4'hb):(1'h0)] wire453;
  reg [(3'h7):(1'h0)] reg452 = (1'h0);
  reg [(5'h12):(1'h0)] reg451 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg450 = (1'h0);
  reg [(5'h12):(1'h0)] reg449 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg448 = (1'h0);
  wire [(4'hc):(1'h0)] wire447;
  wire signed [(2'h3):(1'h0)] wire446;
  wire [(4'hd):(1'h0)] wire445;
  reg signed [(4'h9):(1'h0)] reg444 = (1'h0);
  reg [(3'h7):(1'h0)] reg443 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire442;
  reg signed [(3'h6):(1'h0)] reg441 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg440 = (1'h0);
  reg [(4'hb):(1'h0)] reg439 = (1'h0);
  wire [(3'h4):(1'h0)] wire382;
  wire [(5'h14):(1'h0)] wire383;
  reg [(3'h7):(1'h0)] reg384 = (1'h0);
  reg [(5'h15):(1'h0)] reg385 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg386 = (1'h0);
  reg [(5'h15):(1'h0)] forvar387 = (1'h0);
  reg [(5'h13):(1'h0)] reg388 = (1'h0);
  reg [(5'h15):(1'h0)] reg389 = (1'h0);
  reg [(3'h4):(1'h0)] reg390 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg391 = (1'h0);
  reg [(3'h5):(1'h0)] reg392 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg393 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg394 = (1'h0);
  reg [(5'h10):(1'h0)] reg395 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire396;
  wire [(5'h13):(1'h0)] wire397;
  wire signed [(5'h11):(1'h0)] wire398;
  wire [(5'h15):(1'h0)] wire437;
  assign y = {wire535,
                 wire455,
                 wire454,
                 wire453,
                 reg452,
                 reg451,
                 reg450,
                 reg449,
                 reg448,
                 wire447,
                 wire446,
                 wire445,
                 reg444,
                 reg443,
                 wire442,
                 reg441,
                 reg440,
                 reg439,
                 wire382,
                 wire383,
                 reg384,
                 reg385,
                 reg386,
                 forvar387,
                 reg388,
                 reg389,
                 reg390,
                 reg391,
                 reg392,
                 reg393,
                 reg394,
                 reg395,
                 wire396,
                 wire397,
                 wire398,
                 wire437,
                 (1'h0)};
  assign wire382 = {wire381, (8'hbc)};
  assign wire383 = $unsigned({wire380});
  always
    @(posedge clk) begin
      reg384 = $unsigned(((|(wire380 ?
              (wire382 ? wire379 : wire380) : $signed(wire379))) ?
          $unsigned($signed(wire380[(1'h1):(1'h1)])) : wire380));
      reg385 <= ($unsigned(((((8'h9f) | wire382) ~^ (wire378 ?
              wire381 : (8'hbc))) != (&(~wire383)))) ?
          $signed((((wire383 ? (8'ha5) : (8'h9f)) ?
                  (^wire379) : (wire380 ? (8'h9f) : reg384)) ?
              $signed((|wire382)) : wire380[(1'h0):(1'h0)])) : ((!wire380) ?
              (^~$signed(wire380[(1'h0):(1'h0)])) : {((wire380 ?
                          wire382 : wire380) ?
                      $unsigned(wire379) : (wire378 <= wire381)),
                  $unsigned($signed(wire382))}));
      reg386 <= {reg384[(2'h3):(2'h3)]};
    end
  always
    @(posedge clk) begin
      for (forvar387 = (1'h0); (forvar387 < (1'h0)); forvar387 = (forvar387 + (1'h1)))
        begin
          reg388 <= $signed((!wire381[(3'h5):(2'h3)]));
          reg389 <= $unsigned(($unsigned(wire380) * wire380));
          reg390 <= $signed((((^((8'h9f) + (8'h9f))) && $signed((8'had))) ?
              $unsigned((&(!forvar387))) : ($signed((reg385 <<< reg386)) <<< $signed(((7'h44) <= reg384)))));
          reg391 <= wire378[(3'h4):(2'h2)];
        end
      reg392 = reg385;
      reg393 = {wire382, reg386};
      reg394 <= $unsigned($signed((((reg388 ? wire378 : reg392) << ((8'had) ?
              wire379 : reg391)) ?
          ($unsigned((8'hb7)) != (reg384 ?
              (8'haa) : reg384)) : (reg388[(4'h8):(3'h7)] ?
              (reg392 ? wire379 : reg389) : $unsigned(wire379)))));
      reg395 <= $unsigned(($unsigned((~(wire380 < (8'hb5)))) ?
          $signed((!$signed(wire381))) : $unsigned({wire383})));
    end
  assign wire396 = ($signed((!(8'ha5))) ? reg390[(1'h1):(1'h0)] : (8'ha3));
  assign wire397 = ({($signed(reg388[(4'hf):(3'h4)]) ?
                               $signed({reg384, reg384}) : reg384),
                           $unsigned((forvar387[(3'h4):(2'h3)] || wire383))} ?
                       forvar387[(3'h5):(3'h5)] : ($signed(reg392[(3'h4):(2'h2)]) ?
                           (~^wire381) : (reg391[(4'h8):(3'h6)] ?
                               (+{reg390, wire382}) : $signed({wire383}))));
  assign wire398 = (&(8'hbc));
  module399 modinst438 (wire437, clk, reg386, wire381, forvar387, reg393, reg390);
  always
    @(posedge clk) begin
      reg439 = $signed({(wire380[(3'h6):(2'h2)] < (8'h9e))});
      reg440 <= (&(reg390[(1'h1):(1'h1)] ?
          {{wire437[(3'h5):(2'h3)]}, ((~|wire380) < (^~wire379))} : wire382));
      reg441 <= reg393[(4'hf):(1'h0)];
    end
  assign wire442 = forvar387[(2'h2):(1'h0)];
  always
    @(posedge clk) begin
      reg443 <= $signed((&(reg394[(1'h1):(1'h0)] & $signed(wire442))));
      reg444 <= $signed((|(8'haa)));
    end
  assign wire445 = $signed({wire396, reg389[(4'hc):(3'h7)]});
  assign wire446 = forvar387[(4'he):(2'h3)];
  assign wire447 = $unsigned({{$signed((reg386 & reg395)),
                           $unsigned((~^wire381))},
                       $unsigned(wire396[(1'h1):(1'h0)])});
  always
    @(posedge clk) begin
      reg448 <= reg389[(5'h12):(4'h8)];
    end
  always
    @(posedge clk) begin
      reg449 <= $unsigned({reg384[(2'h2):(1'h0)],
          (((reg389 >= wire442) ? (8'ha5) : {reg394, wire383}) ?
              $unsigned($signed(wire383)) : reg395)});
      reg450 <= (8'hbb);
      reg451 <= wire446[(2'h3):(2'h3)];
      reg452 <= (&$signed($unsigned(($signed(wire442) ^ (wire437 ?
          wire379 : (8'hac))))));
    end
  assign wire453 = $signed(wire445);
  assign wire454 = $unsigned(((|$signed((reg394 ? (8'h9e) : (8'hab)))) ?
                       $unsigned(((8'hb2) ^~ $signed(reg386))) : ($unsigned((-wire382)) << $signed(reg388[(4'hb):(2'h2)]))));
  assign wire455 = $signed((~wire447[(4'hb):(3'h4)]));
  module456 modinst536 (wire535, clk, forvar387, wire378, reg385, reg439);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module456  (y, clk, wire460, wire459, wire458, wire457);
  output wire [(32'h1ba):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire460;
  input wire signed [(5'h15):(1'h0)] wire459;
  input wire signed [(5'h15):(1'h0)] wire458;
  input wire signed [(4'hb):(1'h0)] wire457;
  reg signed [(5'h13):(1'h0)] reg534 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg533 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg532 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg531 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar529 = (1'h0);
  reg [(2'h3):(1'h0)] forvar526 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg530 = (1'h0);
  reg [(3'h7):(1'h0)] reg529 = (1'h0);
  reg [(2'h3):(1'h0)] reg528 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg527 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg526 = (1'h0);
  reg [(4'ha):(1'h0)] reg525 = (1'h0);
  reg [(4'h9):(1'h0)] reg524 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg523 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg522 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar521 = (1'h0);
  reg [(4'h8):(1'h0)] reg520 = (1'h0);
  reg [(5'h13):(1'h0)] reg519 = (1'h0);
  reg [(2'h3):(1'h0)] forvar518 = (1'h0);
  reg [(5'h13):(1'h0)] reg517 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire516;
  wire [(4'hf):(1'h0)] wire515;
  reg signed [(4'he):(1'h0)] reg514 = (1'h0);
  reg [(3'h5):(1'h0)] reg513 = (1'h0);
  reg [(4'h9):(1'h0)] reg512 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire510;
  reg [(5'h13):(1'h0)] reg469 = (1'h0);
  reg [(5'h15):(1'h0)] reg468 = (1'h0);
  reg [(5'h14):(1'h0)] reg467 = (1'h0);
  reg [(5'h14):(1'h0)] reg466 = (1'h0);
  reg [(4'h8):(1'h0)] reg465 = (1'h0);
  wire [(5'h15):(1'h0)] wire464;
  wire signed [(5'h11):(1'h0)] wire463;
  wire [(4'h9):(1'h0)] wire462;
  wire [(4'hd):(1'h0)] wire461;
  assign y = {reg534,
                 reg533,
                 reg532,
                 reg531,
                 forvar529,
                 forvar526,
                 reg530,
                 reg529,
                 reg528,
                 reg527,
                 reg526,
                 reg525,
                 reg524,
                 reg523,
                 reg522,
                 forvar521,
                 reg520,
                 reg519,
                 forvar518,
                 reg517,
                 wire516,
                 wire515,
                 reg514,
                 reg513,
                 reg512,
                 wire510,
                 reg469,
                 reg468,
                 reg467,
                 reg466,
                 reg465,
                 wire464,
                 wire463,
                 wire462,
                 wire461,
                 (1'h0)};
  assign wire461 = {$signed($signed($signed(wire457))), wire460[(4'he):(3'h4)]};
  assign wire462 = $signed($signed((wire458 || wire460[(3'h4):(1'h0)])));
  assign wire463 = ($signed({(~&wire459[(3'h7):(2'h3)])}) + wire461);
  assign wire464 = wire459;
  always
    @(posedge clk) begin
      reg465 <= (8'h9e);
      reg466 <= ($unsigned((wire462[(3'h5):(2'h2)] >= reg465)) - reg465);
      reg467 <= wire459[(4'hc):(3'h4)];
      reg468 <= wire459;
      reg469 = ($signed($unsigned($signed($unsigned(wire463)))) < ((($signed(reg465) * $unsigned(wire461)) ?
          (wire461[(4'h9):(4'h9)] ?
              wire464[(4'h8):(3'h6)] : (wire457 ~^ (7'h40))) : wire463[(2'h3):(2'h3)]) + wire459));
    end
  module470 modinst511 (.wire471(reg469), .y(wire510), .clk(clk), .wire472(wire459), .wire473(wire463), .wire474(reg467));
  always
    @(posedge clk) begin
      reg512 <= $unsigned(($unsigned(reg469) != $signed(wire510)));
      reg513 <= reg466;
      reg514 <= wire464[(5'h12):(4'he)];
    end
  assign wire515 = wire460[(3'h4):(1'h1)];
  assign wire516 = reg513;
  always
    @(posedge clk) begin
      reg517 <= wire510;
      for (forvar518 = (1'h0); (forvar518 < (3'h4)); forvar518 = (forvar518 + (1'h1)))
        begin
          reg519 = (&wire515[(4'h8):(3'h6)]);
          reg520 <= (wire458 ? wire516[(2'h3):(1'h0)] : $signed(reg517));
          for (forvar521 = (1'h0); (forvar521 < (1'h0)); forvar521 = (forvar521 + (1'h1)))
            begin
              reg522 = wire463;
            end
          reg523 <= $signed($unsigned((reg513 - forvar521[(5'h15):(2'h3)])));
          reg524 <= wire510[(4'hb):(2'h3)];
        end
      reg525 <= $signed((reg519[(4'h8):(3'h7)] << reg519[(4'hd):(4'hc)]));
      if (((forvar521[(2'h3):(1'h1)] ?
          (forvar521 < (reg512 >>> forvar521[(4'h9):(2'h3)])) : wire457[(3'h4):(3'h4)]) > (|(~reg465))))
        begin
          reg526 <= wire510;
          reg527 <= wire460[(3'h4):(1'h0)];
          reg528 = wire459;
          reg529 <= ((((7'h43) < (~^wire460)) * (-reg517)) >> (wire515 ?
              (((8'hbe) ? (wire457 * wire463) : wire464) ?
                  wire516 : wire464) : $signed({$unsigned((8'hba)),
                  (^~(7'h44))})));
          reg530 <= (reg520 ~^ reg519[(5'h13):(1'h0)]);
        end
      else
        begin
          for (forvar526 = (1'h0); (forvar526 < (2'h2)); forvar526 = (forvar526 + (1'h1)))
            begin
              reg527 <= (+(^~(~^(reg468[(5'h10):(3'h5)] ?
                  reg469[(4'h8):(3'h5)] : (reg524 << reg529)))));
              reg528 <= $unsigned((((reg530 ? (reg468 | reg529) : {wire463}) ?
                      ({reg526} & reg468) : $unsigned((^~reg527))) ?
                  reg469 : (^$signed({reg514}))));
            end
          for (forvar529 = (1'h0); (forvar529 < (1'h0)); forvar529 = (forvar529 + (1'h1)))
            begin
              reg530 <= wire458[(3'h7):(1'h1)];
            end
          reg531 = $unsigned({forvar521,
              ($signed($unsigned(reg529)) > (reg468[(4'he):(3'h6)] <<< reg522[(2'h3):(2'h3)]))});
          reg532 <= wire460;
          reg533 <= ((({reg525, (reg528 ? (8'hbe) : reg529)} ?
                      ({reg528} ?
                          (reg520 ?
                              reg532 : wire462) : reg467[(2'h3):(1'h1)]) : reg517) ?
                  reg527 : wire516) ?
              ((reg532[(4'hb):(1'h0)] ~^ (-(reg531 ? reg524 : wire458))) ?
                  (~$unsigned((&(8'hbf)))) : $signed(((reg517 ?
                      reg532 : wire516) || (reg531 || reg522)))) : $signed({$unsigned((wire458 ~^ reg514)),
                  $unsigned((reg527 ? reg519 : reg530))}));
        end
      reg534 <= $signed((8'haf));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module399
#( parameter param436 = (&{{(8'hbd)}, (~^(((8'hae) ? (8'hab) : (8'haa)) >= ((8'hb5) > (8'h9d))))}) )
(y, clk, wire404, wire403, wire402, wire401, wire400);
  output wire [(32'h169):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire404;
  input wire [(4'h8):(1'h0)] wire403;
  input wire [(5'h12):(1'h0)] wire402;
  input wire [(4'hf):(1'h0)] wire401;
  input wire signed [(2'h2):(1'h0)] wire400;
  reg signed [(5'h13):(1'h0)] reg435 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg434 = (1'h0);
  reg [(3'h5):(1'h0)] reg433 = (1'h0);
  reg [(4'he):(1'h0)] reg432 = (1'h0);
  reg [(4'h9):(1'h0)] reg431 = (1'h0);
  reg [(4'h9):(1'h0)] forvar430 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar429 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg428 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg427 = (1'h0);
  reg [(3'h7):(1'h0)] reg426 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg425 = (1'h0);
  reg [(4'h8):(1'h0)] reg424 = (1'h0);
  reg [(4'hb):(1'h0)] reg423 = (1'h0);
  reg [(3'h6):(1'h0)] reg422 = (1'h0);
  wire [(4'h9):(1'h0)] wire421;
  reg signed [(4'he):(1'h0)] reg420 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg419 = (1'h0);
  reg [(3'h4):(1'h0)] reg418 = (1'h0);
  reg signed [(4'he):(1'h0)] reg417 = (1'h0);
  reg [(5'h12):(1'h0)] reg416 = (1'h0);
  reg [(3'h5):(1'h0)] reg415 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg414 = (1'h0);
  reg [(5'h12):(1'h0)] reg413 = (1'h0);
  reg [(5'h13):(1'h0)] reg412 = (1'h0);
  reg [(2'h3):(1'h0)] reg411 = (1'h0);
  reg [(5'h15):(1'h0)] reg410 = (1'h0);
  reg [(5'h12):(1'h0)] reg409 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg408 = (1'h0);
  reg [(4'ha):(1'h0)] reg407 = (1'h0);
  reg [(5'h10):(1'h0)] reg406 = (1'h0);
  reg [(3'h7):(1'h0)] reg405 = (1'h0);
  assign y = {reg435,
                 reg434,
                 reg433,
                 reg432,
                 reg431,
                 forvar430,
                 forvar429,
                 reg428,
                 reg427,
                 reg426,
                 reg425,
                 reg424,
                 reg423,
                 reg422,
                 wire421,
                 reg420,
                 reg419,
                 reg418,
                 reg417,
                 reg416,
                 reg415,
                 reg414,
                 reg413,
                 reg412,
                 reg411,
                 reg410,
                 reg409,
                 reg408,
                 reg407,
                 reg406,
                 reg405,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg405 <= ((-$signed(((wire403 ? wire402 : wire401) ?
              {wire400} : wire403[(1'h0):(1'h0)]))) ?
          $signed(wire400) : $signed($signed((wire400[(1'h1):(1'h1)] ^~ wire402[(4'ha):(2'h3)]))));
      reg406 <= ((~&((~&wire404) << ((!wire404) * wire400[(1'h0):(1'h0)]))) || (wire400[(2'h2):(1'h0)] ?
          wire403 : $signed({(!wire404)})));
    end
  always
    @(posedge clk) begin
      reg407 <= reg405;
      reg408 <= $unsigned((&({$signed(wire404), wire402[(2'h2):(1'h1)]} ?
          $signed(reg407[(2'h3):(2'h2)]) : $signed($unsigned(reg407)))));
      reg409 <= wire404;
    end
  always
    @(posedge clk) begin
      reg410 <= ($signed($unsigned(reg405)) <<< wire401[(3'h4):(2'h2)]);
      reg411 = reg405[(3'h6):(2'h2)];
    end
  always
    @(posedge clk) begin
      reg412 = reg410;
      reg413 = $unsigned((({wire402[(4'hf):(2'h2)], (wire404 != reg409)} ?
          ((^reg408) ?
              ((8'hbb) ?
                  (8'ha8) : wire404) : $unsigned(reg405)) : (&(wire402 == reg409))) <= (7'h44)));
      reg414 <= reg407;
      reg415 <= $signed(wire401);
    end
  always
    @(posedge clk) begin
      reg416 <= $unsigned({reg411[(2'h3):(2'h2)]});
      reg417 <= {$signed((({reg411} ?
              (reg415 ^ reg407) : {wire400, reg413}) << (8'haf)))};
      reg418 = $unsigned($signed((8'ha4)));
      reg419 <= $unsigned((^~$signed(reg410[(3'h7):(2'h3)])));
    end
  always
    @(posedge clk) begin
      reg420 <= (~&{$signed((^$unsigned(reg413)))});
    end
  assign wire421 = $signed(((($signed(wire401) >>> {wire401}) + {$unsigned((8'ha2))}) ?
                       $signed($signed((reg409 >> (8'ha9)))) : {$signed(wire400[(1'h1):(1'h0)]),
                           reg413[(4'he):(4'hb)]}));
  always
    @(posedge clk) begin
      reg422 <= ($unsigned(((+$unsigned((8'haf))) | ($unsigned(reg408) >= reg409))) ?
          (($unsigned({wire421, (8'hb6)}) ?
                  $unsigned($signed((8'hab))) : (-(reg412 && reg418))) ?
              wire400[(1'h0):(1'h0)] : (reg414[(3'h5):(1'h1)] ?
                  reg410[(1'h1):(1'h0)] : $unsigned((reg408 ?
                      reg410 : wire404)))) : (reg407[(4'h9):(1'h1)] ?
              reg407 : ((~$unsigned(wire402)) ?
                  reg405 : ((wire400 ?
                      (7'h43) : reg405) < (reg406 + (8'hb5))))));
      reg423 <= wire400;
      reg424 <= $signed($unsigned((reg418 ?
          (^~reg423[(4'h8):(3'h5)]) : wire403[(1'h1):(1'h0)])));
    end
  always
    @(posedge clk) begin
      reg425 <= wire400;
      reg426 <= wire403[(2'h3):(1'h0)];
      reg427 <= $signed($signed(reg419[(1'h1):(1'h0)]));
      reg428 <= $signed((|(reg410 || reg425)));
      for (forvar429 = (1'h0); (forvar429 < (2'h2)); forvar429 = (forvar429 + (1'h1)))
        begin
          for (forvar430 = (1'h0); (forvar430 < (2'h3)); forvar430 = (forvar430 + (1'h1)))
            begin
              reg431 <= reg428;
            end
          reg432 = (reg426[(1'h0):(1'h0)] * (-wire402));
          reg433 <= (-$unsigned($signed(reg424[(3'h7):(1'h1)])));
          reg434 <= ($signed((reg424 ? $unsigned((&reg411)) : wire421)) ?
              reg432[(3'h4):(2'h2)] : ($signed({$signed(reg406),
                      reg427[(4'ha):(1'h0)]}) ?
                  (8'hb7) : (((reg426 ?
                      reg416 : reg410) >> reg416) == reg408)));
          reg435 <= reg416[(5'h10):(4'ha)];
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module470
#( parameter param508 = (((-((~(8'hba)) ^ ((8'ha1) ? (8'hb9) : (8'hb0)))) - {(((8'h9d) ~^ (8'h9d)) || {(8'ha4), (7'h44)})}) >>> ({(!(~^(8'ha2)))} ? (((~|(8'hba)) ? (!(8'ha5)) : ((8'hbf) ? (8'hb4) : (8'ha2))) ? (~^((8'h9d) > (8'hb8))) : ((-(8'hbb)) ? {(8'ha9)} : ((8'haa) ? (8'ha9) : (7'h44)))) : {(((8'hb1) || (8'ha8)) ? (|(8'hb8)) : ((8'ha4) - (7'h41))), (^~((8'haa) ^ (8'hbe)))}))
, parameter param509 = param508 )
(y, clk, wire474, wire473, wire472, wire471);
  output wire [(32'h16f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h7):(1'h0)] wire474;
  input wire [(5'h11):(1'h0)] wire473;
  input wire signed [(5'h15):(1'h0)] wire472;
  input wire signed [(5'h13):(1'h0)] wire471;
  wire signed [(5'h10):(1'h0)] wire507;
  reg [(2'h2):(1'h0)] reg506 = (1'h0);
  wire [(3'h6):(1'h0)] wire505;
  wire signed [(4'hf):(1'h0)] wire504;
  wire [(4'hd):(1'h0)] wire503;
  wire [(4'ha):(1'h0)] wire502;
  wire signed [(4'hc):(1'h0)] wire501;
  reg [(4'hc):(1'h0)] reg500 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg499 = (1'h0);
  reg [(5'h13):(1'h0)] reg498 = (1'h0);
  reg [(2'h2):(1'h0)] forvar497 = (1'h0);
  reg [(4'ha):(1'h0)] reg496 = (1'h0);
  reg [(4'he):(1'h0)] reg495 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire494;
  wire [(4'hc):(1'h0)] wire493;
  wire [(5'h15):(1'h0)] wire492;
  reg signed [(5'h11):(1'h0)] reg491 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg490 = (1'h0);
  wire [(4'hd):(1'h0)] wire489;
  reg [(4'h9):(1'h0)] reg488 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg487 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg486 = (1'h0);
  reg [(3'h7):(1'h0)] reg485 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg484 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire483;
  reg signed [(5'h11):(1'h0)] reg482 = (1'h0);
  reg [(2'h2):(1'h0)] reg481 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg480 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg479 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar478 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg477 = (1'h0);
  reg [(5'h12):(1'h0)] reg476 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire475;
  assign y = {wire507,
                 reg506,
                 wire505,
                 wire504,
                 wire503,
                 wire502,
                 wire501,
                 reg500,
                 reg499,
                 reg498,
                 forvar497,
                 reg496,
                 reg495,
                 wire494,
                 wire493,
                 wire492,
                 reg491,
                 reg490,
                 wire489,
                 reg488,
                 reg487,
                 reg486,
                 reg485,
                 reg484,
                 wire483,
                 reg482,
                 reg481,
                 reg480,
                 reg479,
                 forvar478,
                 reg477,
                 reg476,
                 wire475,
                 (1'h0)};
  assign wire475 = ((|wire471) + wire472);
  always
    @(posedge clk) begin
      reg476 <= $unsigned($signed((wire471 + ((wire474 ?
          wire475 : (8'hbb)) < $unsigned(wire474)))));
      reg477 <= (^$unsigned($unsigned({(reg476 > wire472),
          ((8'haa) ^~ (8'had))})));
      for (forvar478 = (1'h0); (forvar478 < (3'h4)); forvar478 = (forvar478 + (1'h1)))
        begin
          reg479 <= {reg476[(4'he):(3'h7)]};
          reg480 <= $signed(wire475);
          reg481 = (^$signed($signed((^~{(8'ha2), (8'hae)}))));
        end
      reg482 <= (|reg477);
    end
  assign wire483 = wire471[(2'h3):(2'h2)];
  always
    @(posedge clk) begin
      reg484 <= $signed(((~({reg481} > reg477)) ?
          wire474[(3'h6):(3'h4)] : (wire483 ~^ ((wire483 ? forvar478 : reg480) ?
              $unsigned(wire474) : wire475))));
      reg485 <= $unsigned(((&(8'hb9)) ?
          wire483 : $unsigned($unsigned(reg481[(2'h2):(1'h1)]))));
      reg486 = $unsigned($signed((~|(!{reg482}))));
      reg487 = $unsigned(({{reg477[(1'h0):(1'h0)], reg486[(2'h2):(1'h1)]}} ?
          wire483 : $signed(((-reg485) ?
              (wire483 ? reg480 : reg476) : reg484))));
      reg488 <= $unsigned($signed(((-reg482[(3'h7):(2'h2)]) >= (((8'haa) ?
          wire473 : reg482) ^ (reg477 ^~ reg479)))));
    end
  assign wire489 = (($signed($unsigned(((7'h42) >>> reg488))) ?
                           (~&reg477) : reg479) ?
                       $signed((|$unsigned((reg486 ?
                           wire471 : reg484)))) : $unsigned(wire471));
  always
    @(posedge clk) begin
      reg490 <= (+reg481);
      reg491 <= $unsigned(wire483);
    end
  assign wire492 = (~|({reg487[(4'h9):(4'h8)],
                           (((8'haa) ? reg477 : reg485) ?
                               ((8'haf) >> reg485) : reg481)} ?
                       (~&reg476) : reg488[(2'h3):(1'h1)]));
  assign wire493 = ($unsigned($unsigned((reg486[(4'ha):(4'h9)] >= $signed(wire474)))) | (!$signed(($unsigned(reg479) ?
                       wire471[(4'hc):(4'hc)] : {reg477}))));
  assign wire494 = reg477[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      reg495 <= wire489[(3'h4):(2'h2)];
      reg496 = wire493;
      for (forvar497 = (1'h0); (forvar497 < (3'h4)); forvar497 = (forvar497 + (1'h1)))
        begin
          reg498 <= (~(!(reg486 + reg479[(4'h9):(3'h7)])));
        end
    end
  always
    @(posedge clk) begin
      reg499 <= ($unsigned($unsigned(({reg488, wire474} ?
          $unsigned(reg496) : $unsigned(reg487)))) - wire489);
      reg500 <= reg495[(4'hc):(4'hc)];
    end
  assign wire501 = reg487[(4'hd):(3'h4)];
  assign wire502 = forvar497;
  assign wire503 = (reg481 + ($unsigned(reg485) == (($signed(reg481) ?
                       (wire492 ^~ (8'hb6)) : ((7'h43) ^~ wire492)) == ((wire501 ?
                           reg481 : reg498) ?
                       (-reg481) : $unsigned(reg481)))));
  assign wire504 = (|(~&{(^~(reg491 ? reg486 : reg495))}));
  assign wire505 = (((^(-(~&reg482))) == (reg500 ?
                           (forvar478 ?
                               $signed(wire493) : $unsigned((8'hb8))) : (~|$unsigned((8'hb1))))) ?
                       (^~reg481) : {reg481[(1'h1):(1'h0)]});
  always
    @(posedge clk) begin
      reg506 <= $unsigned($unsigned($unsigned(reg498[(5'h11):(4'hf)])));
    end
  assign wire507 = reg488;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module647  (y, clk, wire648, wire649, wire650, wire651, wire652);
  output wire [(32'h2b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire648;
  input wire [(5'h13):(1'h0)] wire649;
  input wire signed [(5'h12):(1'h0)] wire650;
  input wire [(4'hc):(1'h0)] wire651;
  input wire signed [(4'hb):(1'h0)] wire652;
  reg signed [(4'hd):(1'h0)] reg799 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire798;
  reg [(5'h12):(1'h0)] reg797 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire795;
  assign y = {reg799, wire798, reg797, wire795, (1'h0)};
  module653 modinst796 (.wire658(wire650), .y(wire795), .wire654(wire651), .clk(clk), .wire657(wire652), .wire656(wire649), .wire655(wire648));
  always
    @(posedge clk) begin
      reg797 <= {wire651[(1'h0):(1'h0)], (~^(8'hac))};
    end
  assign wire798 = (reg797[(4'h8):(2'h3)] & (wire652[(3'h7):(3'h4)] ?
                       $signed((+(reg797 ?
                           wire651 : wire649))) : ($signed(wire648) >= wire651)));
  always
    @(posedge clk) begin
      reg799 <= $signed((~wire650));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module653
#( parameter param794 = ({(((&(8'ha8)) ? (^(8'hae)) : ((7'h42) + (8'hbd))) ? (((8'hbe) ? (8'ha2) : (8'hac)) >> (8'ha9)) : ((|(7'h42)) ? ((8'hbd) ^~ (8'hb3)) : (+(8'h9d))))} ? ((-(((8'hbc) ^~ (8'ha7)) ? ((8'had) == (8'hb5)) : ((8'hb6) || (8'h9e)))) & ((&((8'ha8) * (8'had))) <<< (((8'h9c) ^ (8'ha2)) && ((8'ha2) ? (8'ha2) : (8'ha0))))) : (-((((8'ha3) ? (8'ha2) : (7'h41)) >= ((8'hb4) > (7'h42))) <<< {(~&(8'h9c)), ((8'ha0) ~^ (7'h40))}))) )
(y, clk, wire658, wire657, wire656, wire655, wire654);
  output wire [(32'h23c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h12):(1'h0)] wire658;
  input wire signed [(3'h4):(1'h0)] wire657;
  input wire signed [(5'h13):(1'h0)] wire656;
  input wire [(3'h5):(1'h0)] wire655;
  input wire [(4'hc):(1'h0)] wire654;
  reg [(3'h5):(1'h0)] reg793 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg792 = (1'h0);
  reg [(4'hd):(1'h0)] reg791 = (1'h0);
  reg [(4'h8):(1'h0)] reg790 = (1'h0);
  reg [(2'h3):(1'h0)] reg789 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar788 = (1'h0);
  reg signed [(4'he):(1'h0)] reg787 = (1'h0);
  reg [(5'h13):(1'h0)] reg786 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg785 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg784 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar783 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire782;
  reg [(4'hb):(1'h0)] reg781 = (1'h0);
  reg [(4'ha):(1'h0)] reg780 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg779 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire778;
  reg signed [(4'h9):(1'h0)] reg777 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg776 = (1'h0);
  reg [(2'h2):(1'h0)] reg775 = (1'h0);
  reg [(4'hb):(1'h0)] reg774 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg773 = (1'h0);
  reg [(5'h15):(1'h0)] forvar772 = (1'h0);
  reg [(4'ha):(1'h0)] forvar771 = (1'h0);
  reg [(4'ha):(1'h0)] reg770 = (1'h0);
  reg [(5'h13):(1'h0)] reg769 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg768 = (1'h0);
  wire [(5'h15):(1'h0)] wire766;
  reg [(4'hc):(1'h0)] reg681 = (1'h0);
  reg [(4'he):(1'h0)] reg680 = (1'h0);
  wire [(4'ha):(1'h0)] wire679;
  reg [(3'h7):(1'h0)] reg678 = (1'h0);
  reg [(3'h7):(1'h0)] reg677 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg676 = (1'h0);
  reg [(4'hd):(1'h0)] reg675 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire674;
  wire [(5'h13):(1'h0)] wire673;
  wire [(4'hf):(1'h0)] wire672;
  reg signed [(4'ha):(1'h0)] reg671 = (1'h0);
  reg [(5'h11):(1'h0)] reg670 = (1'h0);
  reg [(4'hb):(1'h0)] forvar669 = (1'h0);
  reg [(3'h7):(1'h0)] reg668 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg667 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg666 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg665 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg664 = (1'h0);
  reg [(4'ha):(1'h0)] forvar663 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg662 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg661 = (1'h0);
  wire [(3'h7):(1'h0)] wire660;
  wire signed [(2'h3):(1'h0)] wire659;
  assign y = {reg793,
                 reg792,
                 reg791,
                 reg790,
                 reg789,
                 forvar788,
                 reg787,
                 reg786,
                 reg785,
                 reg784,
                 forvar783,
                 wire782,
                 reg781,
                 reg780,
                 reg779,
                 wire778,
                 reg777,
                 reg776,
                 reg775,
                 reg774,
                 reg773,
                 forvar772,
                 forvar771,
                 reg770,
                 reg769,
                 reg768,
                 wire766,
                 reg681,
                 reg680,
                 wire679,
                 reg678,
                 reg677,
                 reg676,
                 reg675,
                 wire674,
                 wire673,
                 wire672,
                 reg671,
                 reg670,
                 forvar669,
                 reg668,
                 reg667,
                 reg666,
                 reg665,
                 reg664,
                 forvar663,
                 reg662,
                 reg661,
                 wire660,
                 wire659,
                 (1'h0)};
  assign wire659 = ((-$unsigned($unsigned((&wire655)))) ?
                       $unsigned(($signed($signed(wire654)) ?
                           {$signed(wire654)} : wire658[(3'h4):(1'h1)])) : (^~(+{(!wire654),
                           (8'ha0)})));
  assign wire660 = $unsigned((wire657 >> {$signed((!wire656))}));
  always
    @(posedge clk) begin
      reg661 = ($signed({(((7'h42) ? (8'ha8) : wire658) ~^ ((8'hbf) ?
              wire655 : (8'hbe))),
          (^~wire655[(2'h2):(1'h1)])}) * ((wire660 ?
              wire655[(2'h2):(1'h0)] : (wire658 ?
                  $signed((8'hb5)) : $signed(wire657))) ?
          $unsigned({{wire657},
              {wire656}}) : $signed($unsigned((wire654 + wire655)))));
      reg662 <= (8'haa);
      for (forvar663 = (1'h0); (forvar663 < (1'h0)); forvar663 = (forvar663 + (1'h1)))
        begin
          if ($unsigned((8'hb0)))
            begin
              reg664 <= wire655[(1'h0):(1'h0)];
              reg665 = (((wire655[(2'h3):(1'h1)] == {wire659[(2'h2):(1'h1)],
                      $unsigned(wire658)}) >= wire654) ?
                  wire655 : $signed(wire655[(2'h2):(2'h2)]));
              reg666 <= $signed(reg661);
              reg667 <= (8'h9d);
              reg668 <= reg661[(4'h8):(2'h2)];
            end
          else
            begin
              reg664 <= $signed($unsigned($signed($unsigned($unsigned(reg662)))));
            end
        end
      for (forvar669 = (1'h0); (forvar669 < (2'h2)); forvar669 = (forvar669 + (1'h1)))
        begin
          reg670 <= {forvar669[(2'h2):(1'h0)],
              (reg668[(1'h1):(1'h0)] ?
                  reg664[(4'hf):(4'h8)] : $unsigned({$unsigned(wire654)}))};
        end
      reg671 <= $unsigned((($signed(reg661) ?
              reg665[(2'h2):(1'h0)] : ($unsigned(wire658) + (~|(8'hb0)))) ?
          (reg661[(1'h0):(1'h0)] != (wire657 - {wire654,
              reg667})) : $unsigned(reg668)));
    end
  assign wire672 = ((wire657 ?
                       {(forvar669[(3'h4):(1'h0)] ?
                               {wire658} : reg664[(3'h7):(2'h2)]),
                           (wire654 ?
                               wire658[(4'h9):(1'h1)] : ((8'ha7) > wire655))} : (~&$signed((forvar669 ?
                           reg662 : wire658)))) > (($unsigned((|wire657)) ?
                       wire654 : ((-(8'ha9)) ?
                           reg670[(4'hd):(2'h3)] : $signed(reg664))) >= (~&$unsigned($unsigned((8'hb9))))));
  assign wire673 = $unsigned(reg661);
  assign wire674 = $signed(wire656);
  always
    @(posedge clk) begin
      reg675 = (reg671[(3'h5):(2'h2)] ?
          ((~|$signed($unsigned(wire654))) | reg671[(3'h7):(3'h7)]) : wire655[(1'h1):(1'h0)]);
      reg676 <= ({$unsigned($unsigned({(8'hb5), reg665}))} ?
          (forvar669[(2'h3):(1'h1)] - wire673[(5'h10):(2'h3)]) : (|(wire673 ?
              (!(8'hb4)) : (forvar663 * reg668[(2'h3):(1'h1)]))));
      reg677 <= reg668;
      reg678 <= $unsigned({((~(~|wire658)) ?
              (~(reg677 ? wire660 : reg667)) : $signed((^~reg668))),
          (({(8'hb3)} >>> $unsigned(reg661)) ?
              wire659 : wire658[(3'h7):(1'h1)])});
    end
  assign wire679 = (~$unsigned(reg678[(2'h3):(1'h0)]));
  always
    @(posedge clk) begin
      reg680 <= $signed($signed((~&wire659)));
      reg681 <= (((8'hb4) <<< $signed($signed($signed(reg677)))) ?
          {(((wire660 ? forvar663 : reg666) < (wire660 ? (7'h44) : wire659)) ?
                  forvar663 : reg675[(2'h3):(2'h2)])} : $signed($signed(($unsigned((8'hb9)) ?
              $signed(wire654) : reg670))));
    end
  module682 modinst767 (.clk(clk), .wire685(wire679), .wire683(wire673), .wire686(wire658), .wire684(wire674), .y(wire766));
  always
    @(posedge clk) begin
      reg768 <= ($signed((!wire660)) ?
          reg665[(2'h3):(1'h0)] : forvar669[(4'hb):(3'h7)]);
      reg769 <= (((-(-{reg666, wire658})) + reg681) >= (~&reg671));
      reg770 <= $unsigned((~&{((reg661 ? reg676 : reg680) ?
              $signed((8'hbf)) : $unsigned(wire659)),
          (reg768 > (7'h41))}));
      for (forvar771 = (1'h0); (forvar771 < (1'h1)); forvar771 = (forvar771 + (1'h1)))
        begin
          for (forvar772 = (1'h0); (forvar772 < (2'h3)); forvar772 = (forvar772 + (1'h1)))
            begin
              reg773 = reg769;
              reg774 <= (~&(&reg675));
              reg775 <= (reg768[(1'h0):(1'h0)] << (+(reg681[(4'hb):(4'hb)] ~^ {wire656,
                  wire654})));
            end
          reg776 <= $signed(wire679[(3'h7):(2'h2)]);
          reg777 <= {$signed(((!$unsigned(forvar771)) >= (~|((8'hb3) ^~ forvar669)))),
              ((wire655 + ((wire660 ? reg680 : reg776) <= (reg671 ?
                  (8'hb8) : reg773))) <= wire658)};
        end
    end
  assign wire778 = wire660;
  always
    @(posedge clk) begin
      reg779 <= (wire660 <= $signed(wire778[(3'h7):(2'h2)]));
      reg780 <= reg773[(2'h3):(1'h1)];
      reg781 <= (({reg777[(4'h8):(3'h4)]} && ({(reg671 ? wire658 : (8'had)),
          (reg680 || reg770)} * $unsigned($unsigned(wire659)))) || $signed(reg661[(2'h2):(1'h0)]));
    end
  assign wire782 = reg670[(3'h5):(2'h3)];
  always
    @(posedge clk) begin
      for (forvar783 = (1'h0); (forvar783 < (1'h0)); forvar783 = (forvar783 + (1'h1)))
        begin
          reg784 <= $signed(wire673[(4'hb):(4'h9)]);
          reg785 <= $signed(reg678);
          reg786 = ($signed((~|reg774)) ?
              $unsigned($signed(reg779[(2'h2):(1'h0)])) : reg678);
          reg787 <= ($unsigned($signed(reg664[(4'hc):(2'h2)])) ^ $unsigned(((((8'hb7) * reg779) ?
                  (reg666 >>> reg776) : (+(8'ha1))) ?
              {(wire658 ? (7'h43) : (8'hae))} : (|$signed(reg680)))));
          for (forvar788 = (1'h0); (forvar788 < (2'h3)); forvar788 = (forvar788 + (1'h1)))
            begin
              reg789 <= $unsigned($signed(($unsigned(reg770[(3'h6):(1'h1)]) ^ (wire778 ?
                  {wire674} : reg779))));
              reg790 = ($unsigned($unsigned(reg776[(4'h8):(2'h3)])) ?
                  {(~$signed($signed(reg661))),
                      $unsigned({wire656[(3'h6):(1'h1)]})} : wire655[(2'h2):(1'h1)]);
            end
        end
      reg791 <= reg667[(1'h1):(1'h1)];
      reg792 <= (($signed(reg773[(3'h7):(2'h2)]) ?
              $signed((|$signed((7'h43)))) : (^~(-reg665[(3'h6):(1'h1)]))) ?
          (~&(~^reg677[(1'h0):(1'h0)])) : {$signed(wire778[(4'ha):(1'h0)]),
              reg786[(3'h7):(2'h3)]});
      reg793 <= reg781;
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module682
#( parameter param764 = {(&(~&{((8'haf) ? (8'h9f) : (8'hb7)), (^(8'h9f))}))}
, parameter param765 = ({({(param764 ? param764 : param764)} ? (!{param764}) : (8'hb8)), (!{(param764 ? param764 : param764), (param764 ? (8'ha0) : (8'hb9))})} ? param764 : param764) )
(y, clk, wire683, wire684, wire685, wire686);
  output wire [(32'h92):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h4):(1'h0)] wire683;
  input wire [(4'hb):(1'h0)] wire684;
  input wire signed [(4'ha):(1'h0)] wire685;
  input wire signed [(5'h12):(1'h0)] wire686;
  wire [(3'h5):(1'h0)] wire763;
  reg [(4'hd):(1'h0)] reg762 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg761 = (1'h0);
  reg [(3'h6):(1'h0)] reg760 = (1'h0);
  reg [(5'h11):(1'h0)] reg759 = (1'h0);
  reg [(4'hd):(1'h0)] reg758 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar757 = (1'h0);
  wire [(4'h8):(1'h0)] wire756;
  wire signed [(4'ha):(1'h0)] wire755;
  wire signed [(4'hb):(1'h0)] wire687;
  reg [(5'h13):(1'h0)] reg688 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg689 = (1'h0);
  wire [(4'h9):(1'h0)] wire753;
  assign y = {wire763,
                 reg762,
                 reg761,
                 reg760,
                 reg759,
                 reg758,
                 forvar757,
                 wire756,
                 wire755,
                 wire687,
                 reg688,
                 reg689,
                 wire753,
                 (1'h0)};
  assign wire687 = (($signed((wire686 ? (&(8'hab)) : (-(8'ha7)))) ?
                       (~|{(wire685 <<< wire685),
                           (wire686 ?
                               wire685 : (8'hbe))}) : (8'hac)) ~^ $unsigned((-wire684[(3'h5):(1'h0)])));
  always
    @(posedge clk) begin
      reg688 = (!((~(7'h40)) ?
          $unsigned(wire683[(3'h4):(2'h3)]) : ($unsigned((wire686 ?
              wire683 : (8'hb6))) | (wire684[(1'h1):(1'h1)] < $signed(wire684)))));
      reg689 = wire685[(4'ha):(4'h9)];
    end
  module690 modinst754 (wire753, clk, wire685, wire687, wire686, reg688, wire684);
  assign wire755 = wire686;
  assign wire756 = ((|(~^wire683)) + $unsigned({(!(wire687 && (8'haf)))}));
  always
    @(posedge clk) begin
      for (forvar757 = (1'h0); (forvar757 < (2'h2)); forvar757 = (forvar757 + (1'h1)))
        begin
          reg758 = wire755;
          reg759 = {{wire687[(4'ha):(4'h9)]},
              (~(wire753 & $unsigned($unsigned((8'h9c)))))};
          reg760 <= $signed($unsigned((!(wire686 <= ((8'hbe) ?
              wire684 : wire687)))));
          reg761 <= $signed($unsigned($signed(({wire686,
              wire756} <<< reg758[(3'h5):(1'h1)]))));
          reg762 <= wire684[(2'h3):(2'h2)];
        end
    end
  assign wire763 = wire753[(1'h0):(1'h0)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module690  (y, clk, wire695, wire694, wire693, wire692, wire691);
  output wire [(32'h293):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire695;
  input wire signed [(4'hb):(1'h0)] wire694;
  input wire signed [(5'h12):(1'h0)] wire693;
  input wire signed [(5'h13):(1'h0)] wire692;
  input wire signed [(4'hb):(1'h0)] wire691;
  reg [(5'h10):(1'h0)] reg752 = (1'h0);
  reg [(4'h8):(1'h0)] reg751 = (1'h0);
  reg [(3'h5):(1'h0)] reg750 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg749 = (1'h0);
  reg [(4'hb):(1'h0)] reg748 = (1'h0);
  reg [(2'h3):(1'h0)] forvar747 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg746 = (1'h0);
  reg [(4'ha):(1'h0)] reg745 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg744 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar743 = (1'h0);
  reg [(4'hf):(1'h0)] forvar742 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg741 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg740 = (1'h0);
  reg [(3'h4):(1'h0)] reg739 = (1'h0);
  reg [(5'h12):(1'h0)] reg738 = (1'h0);
  wire [(3'h5):(1'h0)] wire737;
  reg [(5'h10):(1'h0)] reg736 = (1'h0);
  reg [(4'h8):(1'h0)] reg735 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg734 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg733 = (1'h0);
  reg [(4'hf):(1'h0)] forvar732 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar731 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg730 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire729;
  reg signed [(4'hf):(1'h0)] reg728 = (1'h0);
  reg [(2'h3):(1'h0)] reg727 = (1'h0);
  reg [(3'h4):(1'h0)] forvar726 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg725 = (1'h0);
  reg [(4'he):(1'h0)] reg724 = (1'h0);
  reg [(4'ha):(1'h0)] reg723 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar722 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg721 = (1'h0);
  reg signed [(4'he):(1'h0)] reg720 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire719;
  wire [(5'h14):(1'h0)] wire718;
  reg [(5'h13):(1'h0)] reg717 = (1'h0);
  reg signed [(4'he):(1'h0)] reg716 = (1'h0);
  reg [(5'h15):(1'h0)] reg715 = (1'h0);
  reg [(3'h4):(1'h0)] reg714 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar713 = (1'h0);
  reg [(4'h9):(1'h0)] reg712 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar711 = (1'h0);
  reg signed [(4'he):(1'h0)] reg710 = (1'h0);
  reg [(5'h14):(1'h0)] reg709 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg708 = (1'h0);
  wire [(4'hc):(1'h0)] wire707;
  wire signed [(4'he):(1'h0)] wire706;
  reg signed [(4'hc):(1'h0)] reg705 = (1'h0);
  reg [(5'h11):(1'h0)] reg704 = (1'h0);
  reg signed [(4'he):(1'h0)] reg703 = (1'h0);
  reg [(4'hb):(1'h0)] reg702 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg701 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg700 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar699 = (1'h0);
  reg [(2'h2):(1'h0)] reg698 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire697;
  wire signed [(4'ha):(1'h0)] wire696;
  assign y = {reg752,
                 reg751,
                 reg750,
                 reg749,
                 reg748,
                 forvar747,
                 reg746,
                 reg745,
                 reg744,
                 forvar743,
                 forvar742,
                 reg741,
                 reg740,
                 reg739,
                 reg738,
                 wire737,
                 reg736,
                 reg735,
                 reg734,
                 reg733,
                 forvar732,
                 forvar731,
                 reg730,
                 wire729,
                 reg728,
                 reg727,
                 forvar726,
                 reg725,
                 reg724,
                 reg723,
                 forvar722,
                 reg721,
                 reg720,
                 wire719,
                 wire718,
                 reg717,
                 reg716,
                 reg715,
                 reg714,
                 forvar713,
                 reg712,
                 forvar711,
                 reg710,
                 reg709,
                 reg708,
                 wire707,
                 wire706,
                 reg705,
                 reg704,
                 reg703,
                 reg702,
                 reg701,
                 reg700,
                 forvar699,
                 reg698,
                 wire697,
                 wire696,
                 (1'h0)};
  assign wire696 = {wire691[(2'h2):(1'h1)]};
  assign wire697 = wire694;
  always
    @(posedge clk) begin
      reg698 <= $unsigned(wire695);
      for (forvar699 = (1'h0); (forvar699 < (3'h4)); forvar699 = (forvar699 + (1'h1)))
        begin
          reg700 <= $signed($unsigned((((|(8'hbe)) | $signed(wire692)) ?
              ((wire697 >= wire693) == {wire697, wire695}) : forvar699)));
          reg701 <= (wire691[(3'h5):(2'h3)] ?
              ((7'h43) ?
                  (-$unsigned({wire697,
                      wire696})) : wire694) : $signed(wire693));
        end
      reg702 = $unsigned($signed((^~wire696)));
    end
  always
    @(posedge clk) begin
      reg703 <= $signed(reg702);
      reg704 = wire694;
      reg705 = wire694[(4'hb):(3'h6)];
    end
  assign wire706 = wire691;
  assign wire707 = reg703[(2'h3):(1'h0)];
  always
    @(posedge clk) begin
      reg708 <= $unsigned(wire692);
      reg709 = (wire707 ?
          $unsigned($unsigned((~&(reg705 && reg703)))) : $unsigned(wire691[(4'hb):(1'h1)]));
      reg710 <= (wire692 >= ($signed(wire695) || wire695[(3'h6):(3'h4)]));
      for (forvar711 = (1'h0); (forvar711 < (2'h3)); forvar711 = (forvar711 + (1'h1)))
        begin
          reg712 <= (($unsigned($unsigned(reg702)) ?
              $unsigned(($signed((8'hb9)) < (forvar699 >> reg710))) : (((!wire694) < (reg701 << wire697)) && (wire707[(2'h2):(1'h1)] * {reg703,
                  (8'ha1)}))) - (^wire696));
          for (forvar713 = (1'h0); (forvar713 < (1'h0)); forvar713 = (forvar713 + (1'h1)))
            begin
              reg714 <= {(^~(~^(~|$signed(reg703))))};
              reg715 <= wire692;
              reg716 = wire706[(4'he):(4'h8)];
              reg717 <= $signed($unsigned($unsigned(($signed(reg700) && {reg709}))));
            end
        end
    end
  assign wire718 = $signed((~&forvar713[(4'h8):(1'h1)]));
  assign wire719 = (!(|(($signed(reg717) * $unsigned((8'hbc))) ?
                       ({wire693, reg704} ?
                           (~reg698) : (wire694 != (8'hab))) : (&wire691))));
  always
    @(posedge clk) begin
      reg720 = reg709[(4'he):(4'hd)];
      reg721 <= ({(reg714 ? reg720[(4'h9):(2'h3)] : {$unsigned(wire696)}),
              $signed($signed(((7'h44) != reg703)))} ?
          {(^~$signed((reg715 != wire707)))} : $unsigned((($signed(reg709) ?
              wire691[(4'ha):(4'h9)] : forvar699) ^~ (wire696 >>> (!wire695)))));
      for (forvar722 = (1'h0); (forvar722 < (1'h0)); forvar722 = (forvar722 + (1'h1)))
        begin
          reg723 <= $unsigned($signed($signed($signed(reg717))));
          reg724 <= wire718;
          reg725 <= (|reg723);
          for (forvar726 = (1'h0); (forvar726 < (2'h2)); forvar726 = (forvar726 + (1'h1)))
            begin
              reg727 = (8'hb0);
              reg728 <= wire706;
            end
        end
    end
  assign wire729 = ({{(reg698[(1'h1):(1'h0)] ? reg710 : wire695)}} ?
                       ((($signed(reg698) >> reg720[(1'h1):(1'h0)]) ?
                           ((reg698 ? reg727 : reg698) ?
                               reg720[(4'hd):(3'h5)] : $unsigned(reg721)) : (~^(wire696 >> reg698))) || $signed($unsigned(forvar713[(4'he):(4'h8)]))) : (reg705[(4'ha):(3'h6)] ?
                           $unsigned(((reg724 & (7'h40)) || (8'h9d))) : (reg724 ?
                               $unsigned(reg710[(2'h3):(2'h2)]) : {$signed(wire706)})));
  always
    @(posedge clk) begin
      reg730 <= {forvar699};
      for (forvar731 = (1'h0); (forvar731 < (2'h3)); forvar731 = (forvar731 + (1'h1)))
        begin
          for (forvar732 = (1'h0); (forvar732 < (1'h1)); forvar732 = (forvar732 + (1'h1)))
            begin
              reg733 <= forvar731[(4'hd):(2'h3)];
              reg734 = (reg703 ~^ $unsigned({(&((8'had) ?
                      reg733 : forvar722))}));
              reg735 <= wire697[(1'h1):(1'h0)];
              reg736 = ({($unsigned((reg723 ? reg712 : wire729)) ?
                      (~&(^~(8'hbb))) : $signed((~^(8'hb2)))),
                  $signed({(forvar731 << reg704),
                      ((8'hbf) ? wire706 : (8'ha0))})} && (&(((~&wire707) ?
                  $signed(reg730) : $signed(reg728)) != ((wire694 ?
                      reg700 : forvar722) ?
                  (reg702 + wire695) : (reg702 >> reg714)))));
            end
        end
    end
  assign wire737 = $unsigned(reg725[(3'h7):(3'h7)]);
  always
    @(posedge clk) begin
      reg738 <= (+$signed((8'hb0)));
      reg739 <= $unsigned($signed($signed($signed($unsigned(reg730)))));
    end
  always
    @(posedge clk) begin
      reg740 <= wire718[(4'hb):(4'h9)];
      reg741 = (reg735[(3'h5):(2'h3)] | $unsigned((-(^(reg705 ~^ reg740)))));
      for (forvar742 = (1'h0); (forvar742 < (3'h4)); forvar742 = (forvar742 + (1'h1)))
        begin
          for (forvar743 = (1'h0); (forvar743 < (3'h4)); forvar743 = (forvar743 + (1'h1)))
            begin
              reg744 <= (7'h42);
              reg745 <= ($unsigned((!(~^$unsigned(reg721)))) && forvar742[(3'h6):(1'h0)]);
            end
          reg746 <= (reg709[(5'h14):(4'he)] ?
              {((8'h9c) + wire706[(1'h0):(1'h0)]),
                  (forvar711 >= ((wire695 ?
                      reg745 : reg725) + ((8'ha5) <= forvar742)))} : $signed(((forvar722 ?
                  $signed(reg725) : (&reg727)) && ((wire719 ? reg720 : reg698) ?
                  ((7'h43) ? reg698 : reg700) : $unsigned(reg714)))));
          for (forvar747 = (1'h0); (forvar747 < (1'h1)); forvar747 = (forvar747 + (1'h1)))
            begin
              reg748 <= (forvar713[(4'hb):(3'h7)] >> (forvar722[(4'ha):(4'h8)] ?
                  {($unsigned(reg703) == forvar747[(1'h1):(1'h1)]),
                      $unsigned((-reg730))} : (!$unsigned((reg730 * wire696)))));
              reg749 = reg735;
              reg750 <= ($unsigned(((!(forvar742 ? reg702 : wire691)) ?
                  reg727[(2'h3):(1'h1)] : $signed($signed(reg698)))) <<< $signed($signed(($unsigned(reg749) > (^wire697)))));
              reg751 = (^~$signed($unsigned(reg708)));
              reg752 = forvar711[(1'h1):(1'h0)];
            end
        end
    end
endmodule