module top_1
#( parameter param211 = {((&(((8'hb5) ? (8'ha5) : (8'ha6)) ? ((7'h42) ? (8'ha2) : (8'hbd)) : (!(8'hb0)))) == (~({(8'hb3)} ? ((8'hb9) >> (8'ha4)) : ((8'hac) ? (8'hb8) : (8'hbd))))), ({({(8'ha4), (7'h40)} ? ((8'hbd) && (8'ha2)) : ((7'h43) >> (8'h9c)))} ~^ ((((8'ha7) | (8'had)) && ((8'ha1) ? (8'hbb) : (8'ha6))) && ((^(8'h9e)) ? ((8'ha4) >>> (8'hbb)) : (!(8'ha6)))))}
, parameter param212 = param211 )
(y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h225):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire0;
  input wire [(4'hf):(1'h0)] wire1;
  input wire signed [(3'h5):(1'h0)] wire2;
  input wire [(4'ha):(1'h0)] wire3;
  input wire [(4'hd):(1'h0)] wire4;
  reg [(4'hf):(1'h0)] reg210 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg209 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg208 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg207 = (1'h0);
  wire [(4'h8):(1'h0)] wire206;
  wire signed [(4'hb):(1'h0)] wire204;
  wire [(4'hb):(1'h0)] wire203;
  wire signed [(5'h14):(1'h0)] wire202;
  wire signed [(4'he):(1'h0)] wire201;
  wire signed [(5'h13):(1'h0)] wire199;
  wire signed [(5'h12):(1'h0)] wire86;
  reg signed [(4'h8):(1'h0)] reg85 = (1'h0);
  reg [(5'h14):(1'h0)] reg84 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg83 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire82;
  reg signed [(4'hb):(1'h0)] reg5 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg6 = (1'h0);
  reg [(5'h11):(1'h0)] reg7 = (1'h0);
  reg [(4'hc):(1'h0)] reg8 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg9 = (1'h0);
  reg [(5'h12):(1'h0)] reg10 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg11 = (1'h0);
  reg [(4'hf):(1'h0)] reg12 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg13 = (1'h0);
  reg [(2'h2):(1'h0)] reg14 = (1'h0);
  reg [(4'ha):(1'h0)] reg15 = (1'h0);
  reg [(4'hd):(1'h0)] reg16 = (1'h0);
  reg [(4'ha):(1'h0)] reg17 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg18 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg19 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg20 = (1'h0);
  reg [(4'h8):(1'h0)] reg21 = (1'h0);
  reg [(4'ha):(1'h0)] reg22 = (1'h0);
  reg [(4'hf):(1'h0)] reg23 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg24 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg25 = (1'h0);
  reg [(5'h11):(1'h0)] reg26 = (1'h0);
  reg [(3'h4):(1'h0)] reg27 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg28 = (1'h0);
  wire [(5'h13):(1'h0)] wire29;
  wire signed [(4'hb):(1'h0)] wire30;
  wire signed [(3'h6):(1'h0)] wire31;
  wire signed [(5'h10):(1'h0)] wire32;
  wire signed [(5'h15):(1'h0)] wire80;
  assign y = {reg210,
                 reg209,
                 reg208,
                 reg207,
                 wire206,
                 wire204,
                 wire203,
                 wire202,
                 wire201,
                 wire199,
                 wire86,
                 reg85,
                 reg84,
                 reg83,
                 wire82,
                 reg5,
                 reg6,
                 reg7,
                 reg8,
                 reg9,
                 reg10,
                 reg11,
                 reg12,
                 reg13,
                 reg14,
                 reg15,
                 reg16,
                 reg17,
                 reg18,
                 reg19,
                 reg20,
                 reg21,
                 reg22,
                 reg23,
                 reg24,
                 reg25,
                 reg26,
                 reg27,
                 reg28,
                 wire29,
                 wire30,
                 wire31,
                 wire32,
                 wire80,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg5 <= ((+wire1[(2'h2):(1'h0)]) && $unsigned($unsigned($unsigned((8'ha4)))));
      if (({((8'ha5) ?
                  (8'hab) : ((wire3 > wire2) ?
                      ((8'ha9) ? wire4 : reg5) : $signed(wire2)))} ?
          ($signed(((!reg5) ? {wire1, (8'h9e)} : (wire1 ? wire3 : wire2))) ?
              {(wire0[(3'h4):(1'h0)] ?
                      $unsigned(wire4) : (wire2 ?
                          reg5 : wire0))} : wire3[(1'h1):(1'h0)]) : {({(|wire2),
                      (wire4 ? wire0 : wire2)} ?
                  (^~$unsigned(wire1)) : wire1[(1'h0):(1'h0)])}))
        begin
          reg6 <= wire0;
          if ((wire0 << reg6[(1'h1):(1'h0)]))
            begin
              reg7 <= (($unsigned((8'ha7)) ?
                      ($unsigned((wire4 >= wire4)) * $unsigned($signed(wire0))) : (($signed(wire1) * (-wire3)) - (~|(~wire1)))) ?
                  {((!(~^wire0)) ?
                          ((wire0 ^ wire2) <= $unsigned(reg5)) : (~&wire0[(4'h9):(1'h1)]))} : $signed(wire4));
              reg8 <= (+($signed($unsigned((~&reg6))) ?
                  {($unsigned(wire3) ?
                          reg5[(1'h1):(1'h0)] : {wire2,
                              (8'hae)})} : ($unsigned({wire1,
                      wire4}) + (~^$signed(wire3)))));
            end
          else
            begin
              reg7 <= wire2;
              reg8 <= wire0[(2'h3):(1'h0)];
            end
          reg9 <= ((($signed($signed(reg6)) <= ((wire4 || reg5) + {(8'hbc)})) ?
                  (8'ha7) : $unsigned(({wire0, reg5} ?
                      (reg6 || reg5) : (wire4 ? reg7 : reg6)))) ?
              $unsigned($signed(reg6[(3'h6):(2'h2)])) : (reg5[(3'h4):(2'h2)] < (((reg6 && reg7) ?
                      wire2[(1'h0):(1'h0)] : {wire1, wire3}) ?
                  $signed($signed(wire3)) : (reg7 ?
                      $signed(reg5) : $unsigned((7'h42))))));
        end
      else
        begin
          reg6 <= reg5[(1'h1):(1'h0)];
          if ($unsigned((7'h44)))
            begin
              reg7 <= (~^{$signed((wire1 <<< $unsigned((8'haf))))});
              reg8 <= reg7;
            end
          else
            begin
              reg7 <= wire1;
              reg8 <= (reg7[(3'h5):(1'h0)] ?
                  reg6 : ($signed($unsigned(wire4)) != ((~^((8'ha0) * reg8)) <= {{wire3,
                          reg7}})));
              reg9 <= {wire4,
                  (((^~(8'hbe)) ?
                          wire3[(1'h0):(1'h0)] : $signed($unsigned((8'hac)))) ?
                      $signed((+wire2[(3'h4):(1'h1)])) : (~^reg5))};
            end
          reg10 <= {reg5};
          reg11 <= (8'haf);
        end
      reg12 <= reg6[(2'h3):(1'h1)];
      if ($unsigned(({(~(reg11 || reg6)), $unsigned((~^reg9))} ?
          (8'had) : (~((reg9 ? reg11 : wire0) - (~wire4))))))
        begin
          reg13 <= $unsigned($unsigned(wire3[(1'h0):(1'h0)]));
          reg14 <= reg6[(1'h1):(1'h1)];
          reg15 <= wire2;
        end
      else
        begin
          if ($signed(reg15[(4'h8):(3'h6)]))
            begin
              reg13 <= (($signed(reg8[(4'h9):(4'h8)]) ?
                  ((!reg8) ?
                      ({reg12} ^~ (reg10 ?
                          wire2 : wire2)) : $signed((|wire2))) : reg8[(3'h7):(1'h1)]) && $unsigned($signed($unsigned(wire2[(1'h1):(1'h1)]))));
              reg14 <= $unsigned($signed((+((8'ha1) ?
                  reg6 : (reg14 ? wire1 : reg13)))));
              reg15 <= reg12[(3'h4):(2'h2)];
            end
          else
            begin
              reg13 <= (wire1 ? reg10 : $signed(reg11[(3'h5):(2'h3)]));
              reg14 <= (~|reg12);
              reg15 <= reg8[(1'h0):(1'h0)];
              reg16 <= $unsigned(reg5);
              reg17 <= $signed(((wire2 * {(reg12 ? (8'hb5) : wire1)}) ?
                  wire1 : (~|(~&$unsigned(reg6)))));
            end
          if (wire0[(4'he):(4'hc)])
            begin
              reg18 <= (8'hbb);
              reg19 <= reg15;
            end
          else
            begin
              reg18 <= $unsigned(reg6);
              reg19 <= $unsigned(reg11[(1'h0):(1'h0)]);
              reg20 <= ((reg6 ?
                  {($unsigned(reg10) ?
                          $unsigned(reg6) : (reg6 >>> reg18))} : (|(-$signed(wire0)))) * $signed(reg7[(1'h0):(1'h0)]));
              reg21 <= $unsigned(reg17[(3'h4):(3'h4)]);
            end
          reg22 <= ((-reg5[(3'h5):(3'h5)]) ?
              ($signed(($unsigned(reg13) >= (reg14 * reg17))) ?
                  (~|((reg11 < (8'hb7)) ?
                      (~^reg11) : $unsigned(reg16))) : reg21) : (~^{reg14,
                  $unsigned($unsigned(reg18))}));
          reg23 <= reg10[(4'ha):(3'h6)];
          if ((reg16[(2'h3):(2'h3)] >> reg19[(2'h3):(2'h2)]))
            begin
              reg24 <= {{(~&$unsigned((8'ha3))), reg19}};
              reg25 <= $unsigned(((8'ha3) ?
                  reg5[(1'h0):(1'h0)] : (($signed(reg9) < reg11) + (^~$signed(reg22)))));
              reg26 <= $unsigned((wire0[(1'h1):(1'h0)] ?
                  ($unsigned({reg22}) ?
                      wire4[(3'h5):(2'h2)] : $unsigned((reg17 ?
                          (8'hb2) : (8'hb7)))) : reg7));
              reg27 <= reg10;
              reg28 <= reg26[(4'h9):(3'h6)];
            end
          else
            begin
              reg24 <= (((((reg24 >> reg21) * reg28[(1'h0):(1'h0)]) != $unsigned($unsigned(reg11))) ?
                  reg28[(3'h5):(3'h4)] : (8'hb7)) - (reg22[(4'h8):(1'h0)] ?
                  $signed($unsigned(wire3)) : ((((7'h40) ~^ (8'ha9)) >= $unsigned(wire0)) < $signed(reg13))));
              reg25 <= (reg13 ? (reg5 < reg28[(3'h7):(3'h4)]) : wire3);
              reg26 <= reg9;
              reg27 <= $signed(reg5[(3'h5):(2'h2)]);
            end
        end
    end
  assign wire29 = reg9;
  assign wire30 = {($signed($unsigned(reg15)) ?
                          reg17[(1'h1):(1'h1)] : (({reg23} ?
                                  {(7'h41)} : (reg15 ? reg6 : (8'hba))) ?
                              ((&(8'ha5)) ?
                                  {reg13} : {reg18}) : reg6[(3'h6):(2'h2)]))};
  assign wire31 = $signed(reg15[(3'h4):(2'h2)]);
  assign wire32 = $unsigned(wire1[(3'h4):(3'h4)]);
  module33_1 modinst81 (.clk(clk), .wire36(reg25), .y(wire80), .wire38(reg7), .wire37(wire1), .wire35(reg5), .wire34(reg20));
  assign wire82 = (reg15[(1'h1):(1'h0)] & reg18);
  always
    @(posedge clk) begin
      if ($unsigned({$unsigned({$unsigned(reg24), wire4[(3'h4):(1'h1)]})}))
        begin
          reg83 <= (reg25 ?
              $signed((reg21[(3'h4):(1'h0)] ?
                  reg24 : (^~(reg15 ?
                      (7'h42) : reg16)))) : (~^$unsigned(($unsigned(reg10) >>> reg13))));
          reg84 <= $signed(($signed(reg83[(4'h9):(1'h0)]) | {((wire0 | reg12) ?
                  $unsigned(reg15) : $unsigned(reg11)),
              reg23[(2'h3):(2'h3)]}));
        end
      else
        begin
          reg83 <= wire32;
          reg84 <= wire30[(4'h8):(4'h8)];
        end
      reg85 <= wire1;
    end
  assign wire86 = $unsigned((reg11[(1'h0):(1'h0)] >>> ($unsigned(reg15[(3'h4):(2'h3)]) ?
                      ((wire82 | (8'hb0)) == reg84) : reg21)));
  module87_1 modinst200 (.wire90(reg7), .wire88(wire80), .y(wire199), .clk(clk), .wire89(reg10), .wire91(reg19));
  assign wire201 = {((($signed(reg10) ? (reg6 ~^ reg5) : (~&reg23)) ?
                           {reg27[(2'h3):(1'h1)],
                               (wire2 ? reg25 : (7'h41))} : reg9) ^~ reg6),
                       wire80[(5'h13):(4'ha)]};
  assign wire202 = (8'ha4);
  assign wire203 = ((&$signed(reg18[(4'hb):(2'h3)])) || $signed((~^$unsigned($unsigned((8'h9e))))));
  module39_1 modinst205 (.wire41(reg24), .wire43(reg7), .wire42(reg5), .wire40(reg19), .y(wire204), .clk(clk));
  assign wire206 = ((8'had) ? reg21 : (!$unsigned($signed({reg8}))));
  always
    @(posedge clk) begin
      reg207 <= {($signed({$unsigned(wire204)}) ?
              (reg24[(4'h9):(3'h6)] > ((reg28 ?
                  reg26 : wire206) && (~|reg12))) : $signed($unsigned((reg85 ?
                  (8'hb0) : (8'hb0)))))};
      reg208 <= reg207[(1'h1):(1'h0)];
      reg209 <= $signed(wire82[(4'hb):(4'hb)]);
      reg210 <= $unsigned((((~^$signed(wire4)) ?
              $unsigned((^~reg27)) : reg207) ?
          reg11[(1'h1):(1'h0)] : ((wire80[(2'h3):(2'h3)] ?
                  $unsigned(reg14) : (reg23 ? reg15 : (8'hbb))) ?
              $unsigned((reg83 >= (8'hb3))) : reg26)));
    end
endmodule

module module87_1
#( parameter param198 = (^{({(8'haf), ((8'ha1) ? (8'hba) : (8'ha0))} ? (((8'hb5) ? (8'hb1) : (8'hbc)) ? ((8'haa) ~^ (8'hab)) : {(8'ha8)}) : (~&((8'hac) ? (8'ha4) : (8'hb4))))}) )
(y, clk, wire88, wire89, wire90, wire91);
  output wire [(32'hb0):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire88;
  input wire signed [(5'h12):(1'h0)] wire89;
  input wire signed [(5'h11):(1'h0)] wire90;
  input wire [(5'h13):(1'h0)] wire91;
  reg [(4'hc):(1'h0)] reg197 = (1'h0);
  reg [(4'h9):(1'h0)] reg196 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg195 = (1'h0);
  reg [(4'h8):(1'h0)] reg194 = (1'h0);
  reg [(3'h5):(1'h0)] reg193 = (1'h0);
  reg [(4'he):(1'h0)] reg192 = (1'h0);
  reg [(4'hb):(1'h0)] reg191 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg190 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire92;
  wire signed [(3'h4):(1'h0)] wire93;
  wire [(5'h13):(1'h0)] wire148;
  wire [(2'h2):(1'h0)] wire150;
  wire [(3'h7):(1'h0)] wire151;
  wire signed [(4'hf):(1'h0)] wire152;
  reg [(4'h8):(1'h0)] reg153 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg154 = (1'h0);
  wire [(5'h13):(1'h0)] wire188;
  assign y = {reg197,
                 reg196,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 reg191,
                 reg190,
                 wire92,
                 wire93,
                 wire148,
                 wire150,
                 wire151,
                 wire152,
                 reg153,
                 reg154,
                 wire188,
                 (1'h0)};
  assign wire92 = (wire91[(3'h7):(2'h2)] > {(!(wire89[(1'h1):(1'h0)] ?
                          (wire90 ? wire91 : (8'had)) : $unsigned(wire88)))});
  assign wire93 = (wire89[(4'h9):(3'h7)] <= $unsigned($signed({wire92[(3'h4):(2'h2)]})));
  module94_1 modinst149 (wire148, clk, wire91, wire88, wire89, wire90);
  assign wire150 = $unsigned(wire92);
  assign wire151 = (8'hb6);
  assign wire152 = $unsigned($signed($signed({wire92})));
  always
    @(posedge clk) begin
      reg153 <= (~&{((wire88[(3'h4):(2'h3)] >> (^~wire148)) ?
              wire93 : (wire92[(1'h1):(1'h0)] ^~ wire150))});
      reg154 <= wire150[(1'h0):(1'h0)];
    end
  module155_1 modinst189 (wire188, clk, wire151, wire88, wire91, reg153, reg154);
  always
    @(posedge clk) begin
      if ((wire89[(4'h8):(3'h7)] != wire152[(4'h8):(2'h3)]))
        begin
          reg190 <= wire92[(2'h3):(1'h1)];
          reg191 <= $unsigned(({wire148[(4'ha):(2'h3)],
              wire188[(4'hf):(3'h7)]} < ($unsigned((+(8'ha8))) ~^ $unsigned((reg153 ?
              reg154 : reg153)))));
        end
      else
        begin
          reg190 <= (wire151[(1'h0):(1'h0)] ?
              reg154[(1'h1):(1'h1)] : ((&(&((8'hb7) >> wire150))) > ($unsigned({wire91,
                      reg154}) ?
                  reg191 : ($unsigned(wire188) ?
                      (wire150 ? wire90 : wire151) : $signed((8'ha7))))));
          reg191 <= (wire89[(2'h3):(2'h3)] == $signed($unsigned(wire89[(2'h2):(2'h2)])));
          if ((($signed((((8'hbd) ?
              (8'hb9) : wire93) ^ $unsigned((8'haa)))) >>> ($unsigned((^~wire148)) ?
              (^{wire89, wire90}) : (8'hb3))) <<< reg153))
            begin
              reg192 <= (&wire91[(5'h11):(5'h10)]);
            end
          else
            begin
              reg192 <= wire93;
              reg193 <= ((($signed(wire151) ?
                          ($signed(wire151) ? reg191 : reg190) : wire93) ?
                      (~|(((7'h43) ? wire91 : (8'ha7)) ?
                          (reg153 ?
                              wire89 : wire93) : (~|wire151))) : wire148[(1'h0):(1'h0)]) ?
                  $signed((~&$signed(wire188))) : (wire188 <<< wire148));
              reg194 <= $unsigned((-$signed((^~(|wire150)))));
              reg195 <= (~^$signed(((wire188 ?
                  (|(8'had)) : $signed(wire93)) >>> (8'ha8))));
              reg196 <= reg193[(1'h1):(1'h1)];
            end
          reg197 <= wire150;
        end
    end
endmodule

module module33_1
#( parameter param78 = ((~((~{(8'ha7)}) ^~ (~(&(8'hb2))))) ? (((((8'ha6) ? (8'h9d) : (8'hbd)) + {(8'ha9)}) <= {{(8'ha8)}}) ? (((~&(7'h41)) > (+(8'hac))) | (~&(!(8'hb7)))) : (8'hb1)) : (({((8'haf) ? (8'hbc) : (8'ha0))} && ((~^(7'h44)) ? ((7'h44) && (8'hb0)) : ((8'ha6) * (8'hbf)))) >= (({(8'hac)} ? (^~(8'hba)) : {(8'haa), (8'ha6)}) ~^ (~^((8'hbf) ~^ (8'ha1))))))
, parameter param79 = {((|param78) <<< (-param78))} )
(y, clk, wire38, wire37, wire36, wire35, wire34);
  output wire [(32'h92):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hb):(1'h0)] wire38;
  input wire [(4'hf):(1'h0)] wire37;
  input wire signed [(4'hf):(1'h0)] wire36;
  input wire signed [(3'h7):(1'h0)] wire35;
  input wire signed [(5'h15):(1'h0)] wire34;
  wire signed [(3'h4):(1'h0)] wire77;
  wire signed [(5'h11):(1'h0)] wire76;
  reg signed [(4'ha):(1'h0)] reg75 = (1'h0);
  reg [(4'he):(1'h0)] reg74 = (1'h0);
  reg [(5'h10):(1'h0)] reg73 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg72 = (1'h0);
  reg [(3'h5):(1'h0)] reg71 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg70 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg69 = (1'h0);
  wire [(2'h2):(1'h0)] wire68;
  wire [(3'h4):(1'h0)] wire67;
  wire signed [(5'h14):(1'h0)] wire66;
  wire [(2'h3):(1'h0)] wire65;
  wire [(4'he):(1'h0)] wire64;
  wire [(4'hc):(1'h0)] wire62;
  assign y = {wire77,
                 wire76,
                 reg75,
                 reg74,
                 reg73,
                 reg72,
                 reg71,
                 reg70,
                 reg69,
                 wire68,
                 wire67,
                 wire66,
                 wire65,
                 wire64,
                 wire62,
                 (1'h0)};
  module39_1 modinst63 (.clk(clk), .wire41(wire36), .y(wire62), .wire43(wire37), .wire42(wire38), .wire40(wire34));
  assign wire64 = wire62[(3'h7):(3'h4)];
  assign wire65 = {wire36, {wire35}};
  assign wire66 = {wire36[(1'h0):(1'h0)],
                      ({$signed((wire65 ? wire65 : wire65))} ?
                          {wire65,
                              (!((8'hbc) ?
                                  wire38 : (8'hb6)))} : wire36[(2'h2):(2'h2)])};
  assign wire67 = $unsigned(wire36);
  assign wire68 = ((-wire66[(4'ha):(4'h9)]) ?
                      $unsigned((!wire34)) : $unsigned((+(~|wire35[(1'h0):(1'h0)]))));
  always
    @(posedge clk) begin
      reg69 <= ($signed((((wire38 == wire37) ? (-wire36) : {wire66, wire65}) ?
          (wire34 ?
              (wire37 ?
                  wire65 : wire37) : (^~wire68)) : {$unsigned(wire35)})) | $signed(wire68));
    end
  always
    @(posedge clk) begin
      if ({wire38[(4'hb):(4'h9)]})
        begin
          if (wire37[(4'he):(2'h3)])
            begin
              reg70 <= ((wire34 >= wire65) ? wire66[(3'h5):(3'h4)] : wire34);
            end
          else
            begin
              reg70 <= $signed((8'hba));
              reg71 <= {(~|wire37)};
              reg72 <= (reg71 ?
                  $unsigned($unsigned((-wire62[(4'h9):(2'h3)]))) : {reg69});
              reg73 <= $unsigned(($unsigned(reg70[(4'h8):(2'h2)]) ?
                  {(wire65[(1'h0):(1'h0)] ?
                          wire35[(3'h5):(1'h0)] : (~reg71))} : wire66[(2'h2):(1'h0)]));
              reg74 <= $signed((~^($signed($signed(wire37)) << reg70[(2'h2):(1'h0)])));
            end
          reg75 <= {{reg70[(2'h3):(1'h0)]}, reg74[(3'h6):(3'h6)]};
        end
      else
        begin
          if ((wire66 ?
              ($unsigned(reg71) == ($signed((reg74 | wire64)) && $unsigned((&wire64)))) : reg75))
            begin
              reg70 <= $signed($unsigned($signed(reg71[(3'h4):(2'h2)])));
              reg71 <= $signed({reg69});
              reg72 <= (!reg71[(2'h3):(1'h1)]);
            end
          else
            begin
              reg70 <= ((wire62[(3'h6):(2'h3)] ?
                      wire66[(4'hb):(4'ha)] : ($unsigned((wire62 ?
                          reg69 : reg74)) != $unsigned(wire34[(5'h10):(4'h8)]))) ?
                  reg74 : (wire37 <<< ((((8'hab) && reg75) <= $signed(wire37)) ?
                      wire66[(4'hb):(3'h4)] : $signed($unsigned(wire68)))));
              reg71 <= wire65;
              reg72 <= $unsigned({$unsigned($signed((wire64 ^ wire35)))});
            end
          reg73 <= $unsigned($signed(wire66[(3'h5):(2'h2)]));
          reg74 <= ((&reg69[(2'h3):(1'h0)]) | {($signed($unsigned(reg73)) <<< reg69)});
        end
    end
  assign wire76 = $signed(wire34[(1'h1):(1'h1)]);
  assign wire77 = wire68;
endmodule

module module39_1
#( parameter param60 = ((({{(7'h44), (8'hb1)}, (^(8'hb7))} ? (((8'h9e) ? (8'hb0) : (8'ha4)) ? ((8'hbf) ^~ (8'ha2)) : ((8'haa) < (8'haf))) : ((&(8'hac)) ? {(8'haf)} : {(8'ha9)})) ? {(^~((8'ha9) ? (8'ha9) : (8'hbd)))} : ((((8'h9e) ? (8'ha1) : (7'h40)) | (~&(8'hbb))) ? (-(^~(8'hab))) : (~|{(8'ha8), (8'ha0)}))) && (({(8'hb8)} ? (+(8'ha4)) : (~((8'hbf) ? (8'hb8) : (8'hb6)))) ? {{(-(8'haa))}} : {(((8'ha8) >> (8'hb8)) * (~&(7'h40)))}))
, parameter param61 = (param60 != (~^(8'ha3))) )
(y, clk, wire43, wire42, wire41, wire40);
  output wire [(32'he3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h2):(1'h0)] wire43;
  input wire [(4'hb):(1'h0)] wire42;
  input wire [(4'hf):(1'h0)] wire41;
  input wire [(4'ha):(1'h0)] wire40;
  wire [(5'h15):(1'h0)] wire59;
  wire [(5'h13):(1'h0)] wire58;
  wire signed [(5'h12):(1'h0)] wire57;
  wire [(4'he):(1'h0)] wire56;
  wire signed [(4'hc):(1'h0)] wire55;
  wire [(4'h8):(1'h0)] wire54;
  wire [(4'hf):(1'h0)] wire53;
  wire [(3'h7):(1'h0)] wire52;
  wire [(5'h12):(1'h0)] wire51;
  wire [(4'hc):(1'h0)] wire50;
  wire signed [(5'h15):(1'h0)] wire49;
  reg signed [(5'h15):(1'h0)] reg48 = (1'h0);
  wire [(4'h9):(1'h0)] wire47;
  wire signed [(4'ha):(1'h0)] wire46;
  wire [(4'h8):(1'h0)] wire45;
  wire [(4'hd):(1'h0)] wire44;
  assign y = {wire59,
                 wire58,
                 wire57,
                 wire56,
                 wire55,
                 wire54,
                 wire53,
                 wire52,
                 wire51,
                 wire50,
                 wire49,
                 reg48,
                 wire47,
                 wire46,
                 wire45,
                 wire44,
                 (1'h0)};
  assign wire44 = ($unsigned(wire42) ? wire41 : (~|wire42[(2'h2):(2'h2)]));
  assign wire45 = wire40;
  assign wire46 = ($signed($unsigned(wire45[(3'h6):(2'h3)])) ?
                      $signed((^(8'hbd))) : $unsigned(wire45[(4'h8):(2'h3)]));
  assign wire47 = (!wire46[(3'h4):(1'h0)]);
  always
    @(posedge clk) begin
      reg48 <= wire46[(3'h7):(3'h6)];
    end
  assign wire49 = wire45;
  assign wire50 = wire40[(3'h7):(2'h3)];
  assign wire51 = (reg48 << (~{wire40}));
  assign wire52 = wire42[(4'ha):(3'h6)];
  assign wire53 = $signed((~&(7'h43)));
  assign wire54 = $signed((&(wire51[(3'h4):(1'h0)] ?
                      wire46[(4'h8):(1'h1)] : wire42)));
  assign wire55 = wire50;
  assign wire56 = $unsigned({wire40[(1'h1):(1'h0)], ((~^(7'h41)) + wire50)});
  assign wire57 = $signed(wire52[(1'h0):(1'h0)]);
  assign wire58 = $unsigned(reg48[(4'hf):(4'h8)]);
  assign wire59 = ((($signed((!wire42)) > $unsigned((wire54 ?
                          wire57 : (8'ha8)))) ?
                      $unsigned((~|$signed(wire47))) : $unsigned(wire55)) > wire41[(4'hc):(1'h0)]);
endmodule

module module155_1
#( parameter param186 = ((({((8'hae) & (8'hac))} >>> {{(7'h40)}}) << ((((8'hb7) << (8'ha6)) >>> ((8'ha7) >>> (8'hbe))) >>> (+(~^(8'ha6))))) == ((^(~|{(8'hba), (8'hb4)})) ? (((+(8'ha7)) - ((8'ha0) <<< (8'ha9))) ? (((8'hb1) ? (8'h9c) : (8'ha4)) ? {(8'ha9)} : (^(8'hbb))) : ((^(8'h9d)) ? ((8'hb8) >>> (8'ha4)) : ((8'hb2) && (7'h40)))) : (&(((8'hb8) ? (8'hb0) : (8'hac)) ? ((8'haa) ? (8'hbf) : (7'h44)) : (-(7'h41))))))
, parameter param187 = param186 )
(y, clk, wire160, wire159, wire158, wire157, wire156);
  output wire [(32'h109):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h4):(1'h0)] wire160;
  input wire [(5'h15):(1'h0)] wire159;
  input wire [(3'h6):(1'h0)] wire158;
  input wire [(4'h8):(1'h0)] wire157;
  input wire [(5'h10):(1'h0)] wire156;
  reg signed [(4'h9):(1'h0)] reg185 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg184 = (1'h0);
  reg [(3'h5):(1'h0)] reg183 = (1'h0);
  reg [(4'hd):(1'h0)] reg182 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg181 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg180 = (1'h0);
  reg [(4'hc):(1'h0)] reg179 = (1'h0);
  reg [(5'h11):(1'h0)] reg178 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg177 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire176;
  wire [(4'hd):(1'h0)] wire175;
  wire signed [(5'h15):(1'h0)] wire174;
  wire signed [(4'hd):(1'h0)] wire173;
  wire [(4'h8):(1'h0)] wire172;
  wire [(2'h2):(1'h0)] wire171;
  wire [(4'he):(1'h0)] wire170;
  wire [(4'hc):(1'h0)] wire169;
  wire [(4'hb):(1'h0)] wire168;
  wire [(4'he):(1'h0)] wire167;
  wire [(3'h5):(1'h0)] wire166;
  wire signed [(4'h8):(1'h0)] wire165;
  wire signed [(4'ha):(1'h0)] wire164;
  wire [(3'h6):(1'h0)] wire163;
  wire signed [(3'h5):(1'h0)] wire162;
  wire [(4'ha):(1'h0)] wire161;
  assign y = {reg185,
                 reg184,
                 reg183,
                 reg182,
                 reg181,
                 reg180,
                 reg179,
                 reg178,
                 reg177,
                 wire176,
                 wire175,
                 wire174,
                 wire173,
                 wire172,
                 wire171,
                 wire170,
                 wire169,
                 wire168,
                 wire167,
                 wire166,
                 wire165,
                 wire164,
                 wire163,
                 wire162,
                 wire161,
                 (1'h0)};
  assign wire161 = {(~&(~&(^wire158)))};
  assign wire162 = {((wire156[(4'hf):(3'h4)] ?
                               (^~(~&wire158)) : (~|(wire156 ?
                                   wire158 : wire160))) ?
                           (wire158 >> (-wire156)) : (wire159[(4'h8):(1'h1)] ?
                               $signed((~^wire159)) : (~|(+wire161)))),
                       ({$signed(wire161[(3'h7):(2'h3)]),
                           $unsigned({wire156,
                               wire158})} ^ $unsigned((8'hb1)))};
  assign wire163 = ({wire161} ?
                       wire158 : (~^{$signed(wire161),
                           $unsigned(((8'h9f) ? wire160 : wire158))}));
  assign wire164 = (($signed((wire156[(4'hd):(4'hb)] != $unsigned(wire159))) - ((^$signed(wire162)) >> wire156)) >= $signed(($unsigned($unsigned(wire158)) ?
                       wire162 : wire163[(3'h6):(1'h0)])));
  assign wire165 = wire159;
  assign wire166 = (~wire162[(3'h4):(2'h2)]);
  assign wire167 = ($signed(wire158) <<< wire160);
  assign wire168 = wire160[(1'h1):(1'h1)];
  assign wire169 = ($unsigned((8'hae)) ?
                       wire167 : (wire167 ?
                           (wire166[(3'h4):(1'h1)] ^~ wire168[(4'h8):(4'h8)]) : ($signed((^~wire159)) ?
                               ((8'ha0) >>> $unsigned(wire166)) : (~&$signed(wire165)))));
  assign wire170 = {$unsigned($unsigned(wire158)), (!$signed(wire158))};
  assign wire171 = $signed((({(^~wire160), (~|wire167)} ?
                           (wire167[(4'hb):(2'h3)] ?
                               $unsigned(wire170) : $signed(wire158)) : (&wire158)) ?
                       ({wire167[(3'h4):(2'h2)]} && (~&(wire156 ?
                           wire161 : wire156))) : wire160));
  assign wire172 = wire171;
  assign wire173 = $unsigned($signed((((|wire166) ~^ ((8'ha1) ?
                       wire165 : (8'hbe))) + (((8'hbe) ? wire159 : wire172) ?
                       (wire161 >>> wire168) : (~|(8'hb6))))));
  assign wire174 = (!(^wire157[(3'h7):(2'h3)]));
  assign wire175 = $unsigned({($unsigned((7'h43)) >> ((wire174 ?
                               (7'h40) : (8'haf)) ?
                           (wire157 ? wire163 : wire167) : wire168))});
  assign wire176 = wire157;
  always
    @(posedge clk) begin
      if ((&wire170[(3'h5):(1'h1)]))
        begin
          reg177 <= ($signed((8'hb7)) ^ wire172[(3'h4):(2'h2)]);
          if (($unsigned(wire163[(1'h1):(1'h1)]) ?
              ($unsigned($unsigned({wire176})) != (~&$signed({wire162}))) : $signed($unsigned(wire168[(3'h5):(3'h4)]))))
            begin
              reg178 <= ((wire164[(3'h6):(3'h4)] ?
                  (~|$unsigned((8'hbc))) : {{(wire175 + wire172)},
                      wire165[(3'h7):(3'h6)]}) > (7'h42));
              reg179 <= $signed(($signed($signed(wire168[(4'hb):(4'hb)])) && wire175[(3'h6):(2'h3)]));
              reg180 <= (^~$unsigned((&$signed(wire159[(4'hf):(3'h4)]))));
              reg181 <= (-(($unsigned((wire173 ?
                      wire169 : reg179)) ~^ (wire167 ?
                      $unsigned(reg180) : $unsigned((7'h42)))) ?
                  ((|(8'ha5)) ~^ ($unsigned((8'hbf)) >>> wire162[(2'h2):(1'h0)])) : wire175));
            end
          else
            begin
              reg178 <= $signed(wire162);
              reg179 <= {wire157[(1'h1):(1'h0)], $signed(wire168)};
            end
        end
      else
        begin
          if (($unsigned(wire157) ?
              (($signed((wire176 ?
                  wire156 : wire161)) != $signed(wire176[(3'h6):(1'h1)])) <<< (~&((wire176 == wire176) ?
                  (wire158 == wire163) : wire157))) : (wire176[(3'h4):(1'h1)] ?
                  wire171 : $signed(wire170[(4'h8):(3'h7)]))))
            begin
              reg177 <= {(-$signed(wire158))};
            end
          else
            begin
              reg177 <= wire162[(2'h2):(2'h2)];
            end
          reg178 <= $signed((wire175[(3'h5):(1'h1)] ?
              (~|wire175[(4'hb):(2'h3)]) : $unsigned((~&((8'hb1) - wire173)))));
          reg179 <= $signed($unsigned(($signed((wire168 <<< reg181)) <= (~&wire156))));
        end
      reg182 <= ((8'h9e) ? wire165 : $signed(wire160));
      reg183 <= (|(8'ha7));
      reg184 <= wire162[(1'h0):(1'h0)];
      reg185 <= $signed((|wire165));
    end
endmodule

module module94_1
#( parameter param146 = (~|((8'hbd) < (((^~(8'hb8)) > ((8'hb8) ^~ (8'hb1))) >> (((8'hb9) ? (7'h41) : (7'h43)) ? {(7'h42), (8'hb7)} : (&(8'hb1))))))
, parameter param147 = (((~((param146 ? param146 : param146) >= (param146 || param146))) ? param146 : {param146}) ? (8'h9f) : param146) )
(y, clk, wire98, wire97, wire96, wire95);
  output wire [(32'h25d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h2):(1'h0)] wire98;
  input wire signed [(5'h15):(1'h0)] wire97;
  input wire [(3'h5):(1'h0)] wire96;
  input wire signed [(3'h6):(1'h0)] wire95;
  wire [(4'hd):(1'h0)] wire145;
  wire signed [(4'hb):(1'h0)] wire144;
  reg signed [(3'h5):(1'h0)] reg143 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg142 = (1'h0);
  reg [(5'h13):(1'h0)] reg141 = (1'h0);
  reg [(5'h10):(1'h0)] reg140 = (1'h0);
  reg [(4'h9):(1'h0)] reg139 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg138 = (1'h0);
  reg [(4'hf):(1'h0)] reg137 = (1'h0);
  reg [(3'h6):(1'h0)] reg136 = (1'h0);
  reg [(5'h11):(1'h0)] reg135 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg134 = (1'h0);
  reg [(4'h8):(1'h0)] reg133 = (1'h0);
  reg [(5'h10):(1'h0)] reg132 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg131 = (1'h0);
  reg [(5'h15):(1'h0)] reg130 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg129 = (1'h0);
  wire [(5'h12):(1'h0)] wire128;
  wire signed [(4'h8):(1'h0)] wire127;
  wire [(5'h13):(1'h0)] wire126;
  wire signed [(4'hc):(1'h0)] wire125;
  wire [(5'h13):(1'h0)] wire124;
  reg signed [(5'h14):(1'h0)] reg123 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg122 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg121 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg120 = (1'h0);
  reg [(4'h9):(1'h0)] reg119 = (1'h0);
  reg [(2'h3):(1'h0)] reg118 = (1'h0);
  reg [(5'h13):(1'h0)] reg117 = (1'h0);
  reg [(4'hc):(1'h0)] reg116 = (1'h0);
  reg [(3'h4):(1'h0)] reg115 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg114 = (1'h0);
  wire [(3'h6):(1'h0)] wire113;
  wire signed [(5'h11):(1'h0)] wire112;
  wire [(5'h11):(1'h0)] wire111;
  wire [(5'h13):(1'h0)] wire110;
  wire signed [(4'hc):(1'h0)] wire109;
  wire signed [(5'h11):(1'h0)] wire108;
  wire signed [(2'h3):(1'h0)] wire107;
  wire signed [(5'h15):(1'h0)] wire106;
  wire signed [(3'h5):(1'h0)] wire105;
  reg signed [(3'h6):(1'h0)] reg104 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg103 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg102 = (1'h0);
  reg [(4'hb):(1'h0)] reg101 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire100;
  wire signed [(5'h13):(1'h0)] wire99;
  assign y = {wire145,
                 wire144,
                 reg143,
                 reg142,
                 reg141,
                 reg140,
                 reg139,
                 reg138,
                 reg137,
                 reg136,
                 reg135,
                 reg134,
                 reg133,
                 reg132,
                 reg131,
                 reg130,
                 reg129,
                 wire128,
                 wire127,
                 wire126,
                 wire125,
                 wire124,
                 reg123,
                 reg122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 reg117,
                 reg116,
                 reg115,
                 reg114,
                 wire113,
                 wire112,
                 wire111,
                 wire110,
                 wire109,
                 wire108,
                 wire107,
                 wire106,
                 wire105,
                 reg104,
                 reg103,
                 reg102,
                 reg101,
                 wire100,
                 wire99,
                 (1'h0)};
  assign wire99 = wire95;
  assign wire100 = wire97;
  always
    @(posedge clk) begin
      reg101 <= wire99;
      reg102 <= (&(!((~&$unsigned(wire95)) ?
          {(-wire99)} : ((reg101 ? wire98 : wire98) << $unsigned(wire96)))));
      if ($unsigned(((wire95 >> {wire97[(4'h9):(2'h3)]}) ?
          (wire100 ?
              wire100 : {wire96, $signed(wire98)}) : ({reg102[(3'h4):(3'h4)],
                  $unsigned((8'had))} ?
              $signed($signed((8'hb9))) : ($signed(wire99) ?
                  $signed((8'haf)) : reg101[(4'ha):(1'h1)])))))
        begin
          reg103 <= reg102;
        end
      else
        begin
          reg103 <= ((((~|(reg101 ?
              reg102 : wire97)) & reg101) == $unsigned($unsigned($signed(wire96)))) >> (wire99 || reg101[(2'h2):(1'h1)]));
          reg104 <= reg103[(4'h8):(1'h0)];
        end
    end
  assign wire105 = ((reg102 ?
                       reg104[(1'h1):(1'h0)] : $signed((~^$unsigned(wire97)))) && (!(^reg101)));
  assign wire106 = ($unsigned($signed($signed((~wire97)))) & wire95[(3'h5):(2'h2)]);
  assign wire107 = wire96;
  assign wire108 = wire106;
  assign wire109 = ($signed(reg104[(3'h6):(1'h1)]) > ((~&$unsigned($unsigned(wire108))) ?
                       ((+wire95[(3'h4):(1'h0)]) || $signed((~&wire108))) : (!((^wire107) != wire106[(4'ha):(3'h5)]))));
  assign wire110 = $signed($unsigned($unsigned(reg102)));
  assign wire111 = ({wire109[(2'h2):(2'h2)]} ?
                       $unsigned(wire97) : $signed(({((8'hb4) != wire108)} <= {(+reg104),
                           {wire107, wire96}})));
  assign wire112 = wire99;
  assign wire113 = wire98;
  always
    @(posedge clk) begin
      reg114 <= wire113[(3'h5):(3'h4)];
      reg115 <= $signed(((-(+$signed(wire100))) ?
          wire105[(3'h4):(2'h2)] : (&($signed((8'h9e)) ^~ reg104[(2'h2):(2'h2)]))));
      if ($unsigned(((((wire98 && wire109) < {wire105, (8'ha2)}) != wire111) ?
          (({(8'hb4)} ? (wire108 ? reg103 : wire110) : ((8'hba) >= (8'ha1))) ?
              ((^~wire95) >>> (|(8'hb0))) : wire109) : (-wire105[(2'h2):(1'h1)]))))
        begin
          if ((wire110 ?
              wire109 : (~&(((reg101 && reg114) ?
                  (wire108 * reg101) : (!reg114)) | (wire108 ?
                  (-wire112) : ((8'ha9) >>> wire111))))))
            begin
              reg116 <= (-(^~(~((reg115 != (7'h44)) + wire107))));
              reg117 <= {(($signed($signed(wire99)) ?
                          (8'ha4) : $unsigned(reg114)) ?
                      $signed(((wire100 & wire111) ?
                          (wire112 - wire107) : wire107[(1'h1):(1'h0)])) : wire112),
                  (8'ha4)};
              reg118 <= $unsigned(wire109[(4'h8):(3'h6)]);
            end
          else
            begin
              reg116 <= $unsigned(reg116[(4'ha):(4'h8)]);
            end
        end
      else
        begin
          reg116 <= wire105;
          if (reg104[(2'h3):(2'h2)])
            begin
              reg117 <= reg101;
              reg118 <= $signed(({(-wire96),
                  (^(reg118 ? wire105 : wire98))} ~^ wire105[(3'h5):(3'h4)]));
              reg119 <= $signed(reg116[(1'h0):(1'h0)]);
              reg120 <= wire109[(3'h4):(2'h3)];
            end
          else
            begin
              reg117 <= {wire99[(4'hc):(4'hb)],
                  $signed($unsigned($signed((|wire99))))};
              reg118 <= $signed(wire108[(4'ha):(3'h4)]);
              reg119 <= ($signed($signed($signed((wire109 ?
                      reg114 : (7'h43))))) ?
                  (~reg116) : reg117[(5'h13):(4'he)]);
              reg120 <= $unsigned((~^((-(reg120 ?
                  (8'hab) : wire105)) ^ $unsigned((reg117 ?
                  wire109 : wire108)))));
              reg121 <= (+($signed((((8'hb7) - wire98) | (reg120 >> wire99))) >>> {wire100[(1'h1):(1'h0)],
                  ($unsigned(reg118) != reg101)}));
            end
        end
      reg122 <= reg117[(5'h13):(2'h3)];
      reg123 <= $signed(reg120[(4'hf):(4'hf)]);
    end
  assign wire124 = (wire97[(3'h5):(2'h3)] ?
                       ($signed($unsigned(wire110[(5'h10):(4'hc)])) > reg121[(5'h11):(2'h2)]) : ((((wire108 ?
                                   reg115 : wire96) ?
                               (wire111 ?
                                   wire96 : wire110) : $unsigned(wire96)) == wire113) ?
                           ($unsigned(wire113[(2'h2):(2'h2)]) ?
                               wire108[(5'h10):(3'h5)] : $signed($unsigned(reg102))) : ($unsigned($unsigned(wire95)) ?
                               ((reg104 & (8'h9e)) >> {(8'h9c)}) : (~&{(8'ha7),
                                   reg118}))));
  assign wire125 = (reg103[(1'h1):(1'h1)] >= wire111[(3'h4):(1'h1)]);
  assign wire126 = wire113[(3'h5):(3'h5)];
  assign wire127 = $unsigned(wire124[(2'h2):(2'h2)]);
  assign wire128 = {(^(-{reg119[(2'h3):(1'h1)]}))};
  always
    @(posedge clk) begin
      reg129 <= {$signed(($signed(wire112[(4'h9):(3'h7)]) ^ ($unsigned(reg119) ?
              $unsigned(wire112) : wire125)))};
      reg130 <= (wire99[(4'hf):(2'h2)] ?
          {(wire97[(5'h10):(2'h3)] != $signed($signed((8'hb2)))),
              wire96[(2'h3):(1'h1)]} : wire113);
      reg131 <= reg129;
    end
  always
    @(posedge clk) begin
      reg132 <= reg117;
      reg133 <= (reg102 * (~^$signed($unsigned($signed((8'hbf))))));
      reg134 <= {({wire97[(4'h9):(4'h8)]} <<< (~&$unsigned($unsigned((8'hb8))))),
          wire108};
      if (reg114)
        begin
          reg135 <= {reg116[(3'h7):(1'h0)]};
          reg136 <= $signed(($signed(wire111[(4'he):(2'h3)]) << wire112));
          reg137 <= (reg136 > (8'haf));
          reg138 <= $unsigned((wire113[(3'h6):(2'h2)] ?
              (($unsigned(wire100) && wire99) || $signed(wire95[(3'h5):(3'h4)])) : (8'hb1)));
          if ((~($signed((~|(wire110 ~^ reg117))) - {(reg117 | reg131[(2'h3):(2'h2)]),
              (~^{wire108, reg119})})))
            begin
              reg139 <= wire106[(4'he):(4'he)];
              reg140 <= $unsigned($unsigned((8'hb8)));
              reg141 <= wire105[(2'h3):(2'h3)];
            end
          else
            begin
              reg139 <= (($unsigned(reg121[(4'hd):(4'h9)]) ?
                      (wire97[(4'hc):(3'h6)] || ($unsigned(wire100) < (reg140 ?
                          reg121 : (8'hb3)))) : wire125[(4'hb):(1'h1)]) ?
                  {{reg101[(2'h3):(2'h3)]},
                      wire126[(5'h13):(1'h0)]} : (+$signed(((reg115 ?
                          (8'hab) : wire125) ?
                      (reg129 - (8'ha6)) : (~^reg137)))));
              reg140 <= ((&$unsigned((wire100[(1'h0):(1'h0)] ?
                      (~(8'ha4)) : wire96[(1'h1):(1'h1)]))) ?
                  (+((~&(~|reg141)) ?
                      reg118 : {(wire109 ~^ reg101)})) : (wire128 - reg114[(3'h7):(1'h1)]));
              reg141 <= ((8'ha3) || $unsigned((8'hbc)));
              reg142 <= wire105;
            end
        end
      else
        begin
          reg135 <= reg142;
          reg136 <= wire111;
          reg137 <= ($signed(wire109[(3'h5):(2'h3)]) ?
              {{$signed(reg137)}} : (($signed(reg138) ?
                      ($signed(wire127) ?
                          {wire113} : $signed(wire105)) : reg117) ?
                  ($unsigned(((8'ha1) ? wire111 : wire125)) ?
                      reg114[(1'h1):(1'h0)] : (!(wire106 ?
                          wire108 : wire110))) : $signed(((wire126 != reg119) ?
                      (wire96 ? reg103 : reg142) : $unsigned(wire126)))));
          reg138 <= (wire105 ?
              $signed(((8'ha1) ?
                  {wire105,
                      $unsigned(reg116)} : reg104[(3'h6):(1'h1)])) : ((reg131[(4'ha):(3'h6)] ?
                      $unsigned($signed(reg101)) : (|(8'ha2))) ?
                  $unsigned($unsigned((reg118 ?
                      reg103 : reg116))) : $signed((8'hb2))));
        end
      reg143 <= (wire111[(4'hb):(4'ha)] ?
          {reg136,
              $unsigned((+(~|(8'hba))))} : $signed(((8'hb1) ^ $signed((-reg121)))));
    end
  assign wire144 = $signed($signed($signed($unsigned(((8'hae) >= reg139)))));
  assign wire145 = (reg123 ?
                       wire108[(1'h1):(1'h0)] : (&$unsigned({$signed(reg137)})));
endmodule