(* use_dsp48="no" *) (* use_dsp="no" *) module top
#( parameter param140 = (~|(~^(^{(|(7'h40))})))
, parameter param141 = ((~(((param140 ? param140 : param140) ? (^param140) : (~^param140)) && param140)) + param140) )
(y, clk, wire0, wire1, wire2, wire3);
  output wire [(32'h236):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire0;
  input wire [(5'h13):(1'h0)] wire1;
  input wire [(2'h2):(1'h0)] wire2;
  input wire [(4'hd):(1'h0)] wire3;
  wire [(4'hf):(1'h0)] wire139;
  reg [(4'hd):(1'h0)] reg138 = (1'h0);
  reg [(4'ha):(1'h0)] reg137 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg136 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg135 = (1'h0);
  reg [(3'h4):(1'h0)] reg134 = (1'h0);
  reg [(4'he):(1'h0)] reg133 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg132 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg131 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg130 = (1'h0);
  reg signed [(4'he):(1'h0)] reg129 = (1'h0);
  reg [(3'h6):(1'h0)] reg128 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg127 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg126 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire125;
  reg [(4'he):(1'h0)] reg124 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire123;
  wire signed [(4'hb):(1'h0)] wire122;
  reg signed [(5'h15):(1'h0)] reg121 = (1'h0);
  wire [(5'h15):(1'h0)] wire119;
  reg signed [(2'h2):(1'h0)] reg64 = (1'h0);
  reg [(4'h9):(1'h0)] reg63 = (1'h0);
  reg [(2'h3):(1'h0)] reg62 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg61 = (1'h0);
  reg [(4'ha):(1'h0)] reg60 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg59 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg58 = (1'h0);
  reg [(4'hc):(1'h0)] reg57 = (1'h0);
  reg [(4'hb):(1'h0)] reg56 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg55 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg54 = (1'h0);
  wire signed [(4'he):(1'h0)] wire53;
  reg signed [(4'ha):(1'h0)] reg52 = (1'h0);
  reg [(2'h2):(1'h0)] reg51 = (1'h0);
  reg [(3'h7):(1'h0)] reg50 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg49 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg48 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg47 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg46 = (1'h0);
  wire [(5'h14):(1'h0)] wire45;
  wire [(5'h12):(1'h0)] wire44;
  wire signed [(4'hb):(1'h0)] wire43;
  wire [(5'h15):(1'h0)] wire4;
  wire [(5'h12):(1'h0)] wire5;
  wire signed [(5'h14):(1'h0)] wire6;
  wire [(5'h12):(1'h0)] wire41;
  assign y = {wire139,
                 reg138,
                 reg137,
                 reg136,
                 reg135,
                 reg134,
                 reg133,
                 reg132,
                 reg131,
                 reg130,
                 reg129,
                 reg128,
                 reg127,
                 reg126,
                 wire125,
                 reg124,
                 wire123,
                 wire122,
                 reg121,
                 wire119,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 reg55,
                 reg54,
                 wire53,
                 reg52,
                 reg51,
                 reg50,
                 reg49,
                 reg48,
                 reg47,
                 reg46,
                 wire45,
                 wire44,
                 wire43,
                 wire4,
                 wire5,
                 wire6,
                 wire41,
                 (1'h0)};
  assign wire4 = {{(^~wire2[(1'h1):(1'h1)]), (&$signed((^(8'ha4))))}};
  assign wire5 = wire0;
  assign wire6 = (($unsigned((&(~wire1))) > (((8'had) ?
                         wire2 : (wire2 ? wire4 : wire3)) >>> $unsigned({wire1,
                         wire4}))) ?
                     ($unsigned(({wire1} | (8'hbf))) ?
                         ($signed(wire2[(1'h0):(1'h0)]) ?
                             $unsigned(wire4) : $unsigned((+(7'h43)))) : (($unsigned(wire4) ?
                             {wire3} : wire4) ~^ wire5)) : (($signed($signed((8'hb0))) ?
                         (&(wire4 ? wire4 : (8'haf))) : ((~wire2) ?
                             {wire0} : $unsigned(wire2))) || (wire4[(3'h6):(1'h0)] & $unsigned($unsigned((7'h44))))));
  module7 modinst42 (.wire12(wire1), .wire9(wire5), .wire8(wire6), .clk(clk), .y(wire41), .wire11(wire4), .wire10(wire0));
  assign wire43 = (wire0 ?
                      ({$unsigned(wire4[(3'h6):(3'h5)]),
                          ({wire1} ?
                              $signed((8'ha4)) : (8'ha6))} ^ {wire6[(3'h5):(2'h3)],
                          wire6}) : $unsigned($unsigned($signed(wire0))));
  assign wire44 = ({wire0[(3'h4):(2'h2)]} ~^ (wire0[(4'hf):(4'h9)] == $unsigned(($signed(wire6) ?
                      (wire6 ? (8'hb5) : wire5) : $signed((8'hab))))));
  assign wire45 = ({(wire2 ?
                          ((wire41 ? (8'ha0) : wire41) ?
                              $signed(wire41) : ((8'ha1) ?
                                  wire43 : wire5)) : ($signed(wire3) && (wire41 <= wire2))),
                      ((~^$unsigned(wire0)) ?
                          (&(wire5 ?
                              wire43 : wire4)) : $signed($unsigned(wire5)))} || (($signed($unsigned(wire1)) ?
                      $signed($unsigned(wire44)) : {$signed(wire1),
                          wire4[(4'hb):(4'hb)]}) <= wire43[(1'h1):(1'h1)]));
  always
    @(posedge clk) begin
      if ($signed(((+{(wire1 == wire41)}) <= (+$signed(wire0[(3'h5):(1'h0)])))))
        begin
          if ((wire0[(4'hc):(1'h1)] << (((~$unsigned(wire5)) < $unsigned((wire2 & wire43))) & $signed($signed($signed(wire43))))))
            begin
              reg46 <= (|((({wire2} ?
                      wire4[(5'h15):(4'he)] : $unsigned((7'h41))) >> ((^~wire4) ?
                      ((8'ha8) ? wire3 : wire4) : wire1[(5'h13):(3'h4)])) ?
                  ($unsigned(wire41) <= ((~wire2) ?
                      wire5[(4'he):(1'h0)] : {wire0})) : wire2));
            end
          else
            begin
              reg46 <= (~|$unsigned(wire4));
              reg47 <= (8'hba);
              reg48 <= $unsigned(wire2);
            end
          reg49 <= (wire4 ?
              ((((^~wire43) ? $unsigned(reg46) : $signed(wire43)) ?
                      $signed(reg46) : (~^reg46)) ?
                  wire43 : $signed((^~wire5))) : $unsigned((&(8'hbd))));
          reg50 <= $unsigned({(~^(&(wire44 ? wire4 : wire41))),
              $signed($signed($signed((8'h9d))))});
          reg51 <= ((wire1[(1'h0):(1'h0)] ?
              $signed(((wire41 ^ wire0) <= $unsigned((8'hbd)))) : wire6) & ($unsigned((((8'ha8) >= reg47) * wire4)) * $unsigned(reg48)));
        end
      else
        begin
          reg46 <= wire43[(3'h6):(3'h4)];
          reg47 <= $signed({(!(+(^(8'hbf)))), wire43});
          if ($unsigned((wire3[(3'h5):(3'h4)] ?
              (-$unsigned(reg46[(4'hd):(2'h2)])) : $unsigned(reg46[(4'h8):(4'h8)]))))
            begin
              reg48 <= (8'hba);
              reg49 <= wire4;
            end
          else
            begin
              reg48 <= wire1[(5'h11):(1'h1)];
              reg49 <= reg47;
              reg50 <= reg47[(1'h0):(1'h0)];
            end
        end
      reg52 <= ((-$signed(((reg50 ? wire43 : wire6) ?
          (wire0 < reg48) : (^wire3)))) & $signed(reg51));
    end
  assign wire53 = (|reg51);
  always
    @(posedge clk) begin
      reg54 <= reg46;
      if (wire44)
        begin
          reg55 <= wire4[(4'ha):(1'h1)];
          if ($unsigned({$signed((8'ha7)), wire6}))
            begin
              reg56 <= (wire44[(1'h1):(1'h0)] < $signed(($unsigned((~&wire1)) + (reg47 ?
                  (reg51 << (8'hb2)) : (wire5 ? reg47 : (7'h43))))));
              reg57 <= (reg51[(1'h0):(1'h0)] ~^ reg50[(1'h1):(1'h0)]);
              reg58 <= (wire45 || wire43);
            end
          else
            begin
              reg56 <= wire6[(2'h2):(1'h1)];
              reg57 <= reg50;
              reg58 <= reg54[(4'h9):(3'h7)];
            end
          if ({$unsigned($unsigned(reg51))})
            begin
              reg59 <= ((reg51 + {($unsigned(reg58) ~^ reg55[(3'h4):(2'h2)])}) ?
                  $unsigned($signed(((-reg57) & (reg50 <<< (8'had))))) : (wire53[(2'h2):(2'h2)] ?
                      (|(8'hb1)) : $signed(reg52)));
              reg60 <= $unsigned(reg52[(1'h0):(1'h0)]);
              reg61 <= ($unsigned($signed(reg59)) << (~&($unsigned($signed(wire6)) * wire44)));
              reg62 <= ((((wire43[(3'h6):(2'h3)] || (wire1 ?
                      (8'hae) : wire3)) < $unsigned($unsigned(reg49))) ?
                  $unsigned(($signed(reg46) ?
                      (wire44 ?
                          reg60 : wire0) : (~&reg61))) : reg57) && (&(~|{wire41})));
              reg63 <= $signed((wire53 ? reg55 : wire45));
            end
          else
            begin
              reg59 <= (($unsigned(({reg59,
                  reg63} + (^~(8'hbd)))) ^ wire3) >> wire1);
              reg60 <= $signed(wire44);
            end
        end
      else
        begin
          reg55 <= {($signed((((8'ha7) ?
                      (8'ha3) : wire44) ^ wire43[(1'h0):(1'h0)])) ?
                  $signed(((reg63 < wire5) * $signed(wire43))) : $signed(reg48[(4'h9):(3'h4)]))};
          if ($unsigned(wire44))
            begin
              reg56 <= (~&$signed(($signed($unsigned(reg50)) <<< (wire1[(5'h10):(3'h5)] ?
                  wire5[(3'h7):(1'h0)] : reg46[(3'h7):(1'h0)]))));
              reg57 <= $unsigned((|(~$signed((reg57 < reg46)))));
              reg58 <= wire43[(2'h2):(1'h1)];
              reg59 <= $signed((&((-(~^wire4)) ^ ((reg61 ? reg52 : (8'hb0)) ?
                  (reg57 && (8'h9d)) : reg63[(4'h8):(3'h4)]))));
              reg60 <= (~&reg46);
            end
          else
            begin
              reg56 <= reg46;
              reg57 <= $unsigned(({(reg58 ? reg51 : wire3[(4'h8):(3'h7)]),
                  reg59} << $unsigned({{(8'ha9), (8'ha6)}, reg46})));
              reg58 <= $signed($signed(wire0));
            end
          reg61 <= ((|(!$unsigned($signed(reg52)))) >> reg55);
          reg62 <= wire41;
          reg63 <= reg59[(3'h4):(1'h0)];
        end
      reg64 <= ($unsigned(reg54[(4'hd):(2'h2)]) ?
          ((+{wire45[(5'h11):(2'h2)]}) ?
              reg55 : $unsigned($signed(((8'hbc) ?
                  wire53 : wire41)))) : ($signed(reg48[(1'h1):(1'h0)]) ?
              ($unsigned((reg50 ? (8'hbe) : reg52)) ?
                  reg48[(4'h9):(4'h8)] : $unsigned({wire2})) : $signed($signed($unsigned(wire43)))));
    end
  module65 modinst120 (wire119, clk, reg61, wire6, reg60, wire44);
  always
    @(posedge clk) begin
      reg121 <= $signed($signed(($signed(wire5[(5'h12):(5'h10)]) | (reg46 < (!reg46)))));
    end
  assign wire122 = ({reg52[(3'h6):(1'h0)]} < {reg121[(5'h12):(5'h11)],
                       (wire3[(3'h6):(3'h5)] ?
                           wire5 : ($signed(wire44) || $unsigned(reg51)))});
  assign wire123 = ($signed($unsigned($unsigned(reg51[(1'h0):(1'h0)]))) - (wire41[(5'h10):(4'h9)] > $signed({(reg48 ?
                           wire3 : wire6)})));
  always
    @(posedge clk) begin
      reg124 <= reg47[(3'h5):(1'h1)];
    end
  assign wire125 = $signed((8'hb5));
  always
    @(posedge clk) begin
      reg126 <= reg49;
      reg127 <= (8'ha9);
      reg128 <= $unsigned(((&((reg52 ? wire2 : (8'hb3)) ?
              $unsigned(wire3) : reg57[(4'hb):(1'h0)])) ?
          ((-reg52) ~^ wire53) : wire3[(4'ha):(4'ha)]));
      if ((((8'h9f) ?
              ((|((8'hba) ?
                  reg58 : wire0)) <= $signed($unsigned(reg55))) : ((+wire2[(1'h0):(1'h0)]) >= (-reg49[(2'h3):(1'h0)]))) ?
          (($signed((wire53 ?
              wire43 : wire123)) | reg51) | $unsigned(wire125)) : $unsigned(reg59)))
        begin
          reg129 <= reg54;
          reg130 <= ($signed($signed($signed(wire0[(2'h3):(2'h2)]))) ?
              $signed($unsigned($unsigned((reg127 <= wire2)))) : (($unsigned((~|(8'hae))) >>> reg48) ^ wire41[(3'h4):(1'h0)]));
          reg131 <= {reg56, reg61[(4'hb):(4'h8)]};
          reg132 <= (({(|(8'hb0))} ?
                  {(reg61[(4'h9):(4'h9)] ? $unsigned(wire125) : $signed(reg63)),
                      (8'h9c)} : reg48[(4'h9):(3'h6)]) ?
              $unsigned($unsigned(wire122)) : reg58);
        end
      else
        begin
          if ($signed((8'ha8)))
            begin
              reg129 <= $unsigned((((reg55[(1'h1):(1'h0)] ?
                  ((8'haa) ?
                      (8'haf) : wire119) : $signed((8'ha0))) & $signed({reg61})) ^~ reg56[(3'h5):(1'h0)]));
              reg130 <= wire6;
              reg131 <= (~&((reg57 || {$unsigned(reg60)}) + {(+(reg57 ?
                      wire119 : reg64))}));
            end
          else
            begin
              reg129 <= ($unsigned((reg46 << $signed((reg55 | reg129)))) != reg132[(2'h3):(1'h1)]);
              reg130 <= (((~&wire6) ?
                      (^$unsigned((wire1 ?
                          wire43 : wire45))) : reg55[(1'h0):(1'h0)]) ?
                  ($unsigned($unsigned($unsigned((8'ha7)))) >>> (+((reg121 || reg54) & wire0[(4'hd):(3'h5)]))) : reg49);
              reg131 <= ($unsigned((reg64[(2'h2):(2'h2)] * reg48[(1'h0):(1'h0)])) >>> $unsigned(wire45));
            end
          reg132 <= (-$unsigned($unsigned($signed(((8'hb0) > reg126)))));
          if ({$signed(wire0)})
            begin
              reg133 <= reg62[(1'h1):(1'h0)];
              reg134 <= wire4[(3'h7):(1'h0)];
              reg135 <= wire3;
              reg136 <= (|$signed((reg134 ?
                  $signed(reg57) : $unsigned(wire125[(1'h0):(1'h0)]))));
            end
          else
            begin
              reg133 <= reg62;
              reg134 <= (^$unsigned((8'hbb)));
              reg135 <= $unsigned(((+reg133[(4'hc):(2'h2)]) ?
                  ($signed($signed(wire6)) ?
                      (-wire5[(1'h0):(1'h0)]) : $unsigned((+reg129))) : $signed($unsigned(reg128[(3'h6):(1'h0)]))));
              reg136 <= wire41[(4'ha):(2'h2)];
              reg137 <= ($signed($unsigned(wire4[(3'h6):(1'h0)])) ?
                  ((^$signed(wire2)) > (((reg50 ?
                      reg64 : reg57) - (reg48 > reg135)) && wire0[(2'h3):(1'h0)])) : $unsigned({($signed(wire1) - $signed(wire45))}));
            end
        end
      reg138 <= $unsigned(reg137);
    end
  assign wire139 = reg46;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module65
#( parameter param117 = ((+(|((+(8'h9c)) || {(8'hbf)}))) ? ((((~(8'hb1)) ? {(8'ha0), (8'hac)} : ((8'h9f) ? (7'h40) : (8'hb1))) ? (((8'hbf) ? (8'hb7) : (8'hbe)) != ((8'ha2) ? (8'hab) : (8'hb8))) : {(^(8'ha5))}) ? {(((8'hb4) > (8'ha0)) ? {(8'hb9), (8'hb5)} : (~(8'had))), (&(+(8'haa)))} : {({(8'ha8)} ? (|(8'hb9)) : ((8'h9e) ? (7'h44) : (8'ha8))), (~&(~^(8'haa)))}) : (8'ha2))
, parameter param118 = param117 )
(y, clk, wire69, wire68, wire67, wire66);
  output wire [(32'h26f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire69;
  input wire [(5'h14):(1'h0)] wire68;
  input wire [(4'h8):(1'h0)] wire67;
  input wire [(5'h12):(1'h0)] wire66;
  reg [(3'h7):(1'h0)] reg116 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire115;
  wire signed [(4'ha):(1'h0)] wire114;
  wire signed [(4'h9):(1'h0)] wire113;
  wire [(5'h12):(1'h0)] wire112;
  reg signed [(4'hd):(1'h0)] reg111 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg110 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg109 = (1'h0);
  reg [(5'h10):(1'h0)] reg108 = (1'h0);
  wire [(2'h2):(1'h0)] wire107;
  wire [(5'h11):(1'h0)] wire106;
  reg signed [(5'h12):(1'h0)] reg105 = (1'h0);
  reg [(5'h15):(1'h0)] reg104 = (1'h0);
  reg [(3'h7):(1'h0)] reg103 = (1'h0);
  reg [(3'h6):(1'h0)] reg102 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg101 = (1'h0);
  reg [(4'h9):(1'h0)] reg100 = (1'h0);
  reg [(5'h11):(1'h0)] reg99 = (1'h0);
  reg [(5'h11):(1'h0)] reg98 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg97 = (1'h0);
  reg [(4'he):(1'h0)] reg96 = (1'h0);
  reg [(5'h14):(1'h0)] reg95 = (1'h0);
  reg [(4'hc):(1'h0)] reg94 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg93 = (1'h0);
  reg [(5'h10):(1'h0)] reg92 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg91 = (1'h0);
  wire [(4'ha):(1'h0)] wire90;
  wire signed [(3'h7):(1'h0)] wire89;
  wire signed [(5'h15):(1'h0)] wire88;
  wire signed [(4'hb):(1'h0)] wire87;
  wire [(5'h11):(1'h0)] wire86;
  wire signed [(5'h15):(1'h0)] wire85;
  reg signed [(5'h15):(1'h0)] reg84 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg83 = (1'h0);
  reg [(3'h4):(1'h0)] reg82 = (1'h0);
  reg [(4'hf):(1'h0)] reg81 = (1'h0);
  reg [(5'h13):(1'h0)] reg80 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg79 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg78 = (1'h0);
  reg [(3'h7):(1'h0)] reg77 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg76 = (1'h0);
  reg [(4'h8):(1'h0)] reg75 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg74 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire73;
  wire signed [(4'hc):(1'h0)] wire72;
  wire [(4'hd):(1'h0)] wire71;
  wire [(5'h15):(1'h0)] wire70;
  assign y = {reg116,
                 wire115,
                 wire114,
                 wire113,
                 wire112,
                 reg111,
                 reg110,
                 reg109,
                 reg108,
                 wire107,
                 wire106,
                 reg105,
                 reg104,
                 reg103,
                 reg102,
                 reg101,
                 reg100,
                 reg99,
                 reg98,
                 reg97,
                 reg96,
                 reg95,
                 reg94,
                 reg93,
                 reg92,
                 reg91,
                 wire90,
                 wire89,
                 wire88,
                 wire87,
                 wire86,
                 wire85,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 reg80,
                 reg79,
                 reg78,
                 reg77,
                 reg76,
                 reg75,
                 reg74,
                 wire73,
                 wire72,
                 wire71,
                 wire70,
                 (1'h0)};
  assign wire70 = wire69[(1'h0):(1'h0)];
  assign wire71 = $signed(wire68[(5'h10):(4'ha)]);
  assign wire72 = ({wire71} << wire70);
  assign wire73 = wire67;
  always
    @(posedge clk) begin
      if ($unsigned(({{(&wire69), (7'h41)},
          (8'hb5)} || ((+(~|wire68)) && wire71))))
        begin
          if ($signed(wire66[(4'he):(1'h1)]))
            begin
              reg74 <= (8'had);
              reg75 <= reg74[(4'hf):(4'ha)];
              reg76 <= ((reg74 | $unsigned(wire67[(1'h1):(1'h1)])) ?
                  (|$signed((-$signed(reg75)))) : wire69);
              reg77 <= wire73;
              reg78 <= wire70[(2'h2):(1'h0)];
            end
          else
            begin
              reg74 <= wire70;
            end
          reg79 <= (wire67[(1'h1):(1'h1)] >>> $signed(reg74[(2'h3):(1'h1)]));
          reg80 <= $signed(wire66);
          reg81 <= (((((reg75 ? wire72 : (8'hb7)) ?
                  wire66 : wire66) << $unsigned((!reg75))) ?
              ($unsigned((reg75 ? reg78 : wire69)) ?
                  ($signed(wire71) ?
                      (reg78 ?
                          (8'ha1) : (8'haf)) : wire70[(4'h9):(3'h7)]) : $unsigned(reg77[(1'h1):(1'h1)])) : ((wire73 >>> (-(8'hbd))) ?
                  ((reg77 ? wire72 : reg80) ?
                      (reg77 <= wire73) : (!reg80)) : ((reg76 ^ wire71) ?
                      wire72[(4'ha):(3'h7)] : (wire67 ?
                          reg78 : wire67)))) != {$signed((~&reg78)),
              (^~(reg75[(4'h8):(3'h5)] ?
                  $unsigned(reg74) : {wire66, wire72}))});
          reg82 <= (!reg78[(3'h5):(2'h3)]);
        end
      else
        begin
          if (reg76)
            begin
              reg74 <= wire71;
              reg75 <= $unsigned(wire71[(2'h3):(2'h3)]);
              reg76 <= wire73;
              reg77 <= $unsigned($unsigned({reg76}));
              reg78 <= ((^{{reg78[(4'hd):(3'h7)]}}) ?
                  reg80 : reg81[(2'h3):(2'h2)]);
            end
          else
            begin
              reg74 <= (((&$unsigned((wire73 || wire71))) ?
                  ($signed(reg75) ?
                      reg77 : {((8'hb5) ? wire68 : reg80),
                          (reg77 || wire71)}) : wire66[(4'h9):(2'h3)]) == $unsigned($unsigned($signed($signed((8'hae))))));
              reg75 <= reg74[(5'h10):(4'hd)];
              reg76 <= $signed((8'hab));
              reg77 <= $signed({$unsigned((&$signed(wire66)))});
              reg78 <= reg76;
            end
          reg79 <= $unsigned($signed(reg77));
          reg80 <= (8'hb6);
          if (wire73[(4'h8):(3'h5)])
            begin
              reg81 <= ((wire73 >> (+wire68)) ?
                  ((+$unsigned((~^reg81))) | {(reg80 ? (~^reg78) : reg79),
                      $signed((wire70 ?
                          reg82 : wire73))}) : wire71[(3'h5):(1'h1)]);
              reg82 <= wire68[(4'ha):(4'ha)];
              reg83 <= $unsigned(wire70);
              reg84 <= (((((&wire70) ? {reg75} : (reg76 != wire72)) ?
                      (|reg74) : $unsigned(wire72[(2'h3):(1'h0)])) && {{wire69[(4'h8):(2'h3)],
                          reg75},
                      $unsigned((wire69 - wire68))}) ?
                  (reg78[(4'hc):(4'hb)] ?
                      (reg81[(3'h5):(1'h1)] ?
                          reg76[(2'h2):(1'h0)] : $signed((+wire73))) : (wire71[(3'h6):(3'h4)] == (reg81 ?
                          (~&(8'ha5)) : $unsigned(wire69)))) : ($unsigned(((reg81 <= reg75) ?
                          (wire67 ? reg81 : reg74) : reg77[(3'h4):(1'h1)])) ?
                      reg79 : (reg74[(5'h10):(1'h0)] ?
                          wire72[(3'h7):(3'h4)] : (~|$signed(wire69)))));
            end
          else
            begin
              reg81 <= $unsigned($unsigned(((reg78 ?
                      wire72[(1'h1):(1'h1)] : {reg75, wire68}) ?
                  ($signed((8'ha3)) ?
                      (wire66 || reg74) : {reg76, wire69}) : (wire72 ?
                      reg78[(1'h1):(1'h0)] : (reg77 ? reg76 : (7'h41))))));
              reg82 <= reg84[(1'h0):(1'h0)];
            end
        end
    end
  assign wire85 = reg77[(3'h7):(2'h2)];
  assign wire86 = (~&((reg84 ?
                          (reg77[(3'h6):(2'h3)] ?
                              ((8'haf) && wire73) : reg76[(3'h7):(1'h0)]) : $unsigned($signed(wire71))) ?
                      (-{(wire67 ? (8'h9f) : wire70),
                          reg82[(1'h0):(1'h0)]}) : (~(wire72[(4'hb):(3'h4)] ^ $signed((7'h43))))));
  assign wire87 = wire72;
  assign wire88 = ((&(reg83[(2'h3):(1'h0)] ^~ reg81)) ?
                      $unsigned({(~|(-(8'ha5))), reg82}) : (8'ha9));
  assign wire89 = $unsigned((reg78 * wire69[(3'h6):(2'h2)]));
  assign wire90 = reg81;
  always
    @(posedge clk) begin
      reg91 <= (^$unsigned(reg82));
      reg92 <= reg74[(3'h5):(1'h0)];
      if (wire71[(2'h3):(2'h3)])
        begin
          if ($unsigned(((wire68 * $signed(wire67)) ?
              {$signed(reg77[(3'h6):(3'h4)])} : $signed((&(wire89 ?
                  reg77 : (8'h9d)))))))
            begin
              reg93 <= $signed((wire90[(3'h6):(3'h6)] + ((|reg92[(4'h9):(3'h6)]) ?
                  ((reg78 >>> reg76) & {(8'hae)}) : $unsigned($unsigned((8'h9c))))));
              reg94 <= $unsigned($unsigned($signed((&(~^(7'h43))))));
            end
          else
            begin
              reg93 <= $signed((wire71[(2'h3):(2'h2)] ? reg94 : reg74));
              reg94 <= $signed(reg84[(4'hb):(2'h3)]);
              reg95 <= {reg76};
            end
          reg96 <= {$signed(reg93)};
          if (((8'hb6) ?
              $unsigned($unsigned((&$signed(reg93)))) : ({(|reg74[(5'h10):(4'he)]),
                  {(-(8'hbf))}} * wire90)))
            begin
              reg97 <= ((~|((~reg75[(1'h0):(1'h0)]) ?
                      wire67 : ((reg77 ? (8'hb8) : reg95) ?
                          (8'ha1) : wire90[(3'h6):(3'h4)]))) ?
                  ($signed((reg94 + $unsigned((8'hbf)))) ?
                      $unsigned(({(8'hae), reg82} ?
                          wire69 : (~^reg84))) : (~reg79[(3'h5):(3'h4)])) : reg94[(2'h2):(1'h1)]);
            end
          else
            begin
              reg97 <= $signed($unsigned($signed((reg91[(1'h1):(1'h1)] >>> (+reg92)))));
              reg98 <= $unsigned((~wire87[(4'h8):(2'h3)]));
            end
          reg99 <= (&(8'hab));
          if (({wire68} ?
              $unsigned((wire71 ?
                  $unsigned(reg92) : $signed($signed(wire85)))) : (~&(+(wire68[(4'he):(3'h6)] ?
                  wire66 : $unsigned(wire89))))))
            begin
              reg100 <= (wire69 ^~ $unsigned((~|wire72)));
              reg101 <= (($unsigned((&(~^reg81))) ?
                      (8'ha4) : $signed((-$unsigned(reg95)))) ?
                  $signed(reg77[(2'h2):(2'h2)]) : (reg95 || wire71));
              reg102 <= (|$signed(reg80));
              reg103 <= reg100[(2'h2):(1'h0)];
            end
          else
            begin
              reg100 <= $unsigned(reg101);
              reg101 <= $signed((~wire71));
              reg102 <= (~^(reg101[(1'h1):(1'h1)] >= $unsigned({reg83[(1'h1):(1'h0)],
                  (^reg77)})));
              reg103 <= reg101;
            end
        end
      else
        begin
          reg93 <= reg75[(3'h4):(2'h3)];
          reg94 <= (8'h9e);
        end
      reg104 <= $unsigned((|wire89[(1'h0):(1'h0)]));
      reg105 <= reg80;
    end
  assign wire106 = ((reg79 != reg101) ?
                       ($signed((~|$unsigned(reg100))) >= (&(wire89[(3'h4):(2'h2)] < (reg80 <<< (8'h9e))))) : $unsigned((((^reg101) <<< reg102[(2'h2):(2'h2)]) ^ ((reg102 ?
                               reg77 : wire86) ?
                           $unsigned(wire88) : $signed(reg74)))));
  assign wire107 = $unsigned($unsigned(reg84[(3'h6):(1'h1)]));
  always
    @(posedge clk) begin
      reg108 <= reg91;
      reg109 <= $unsigned({reg84[(4'h8):(2'h3)], reg79});
      reg110 <= ((reg77 - ($signed($unsigned((8'hbe))) <= reg77[(1'h0):(1'h0)])) ?
          {reg108[(1'h1):(1'h0)]} : (reg96[(4'ha):(2'h2)] ?
              (^~{wire67}) : (~^$unsigned((reg95 >> reg80)))));
      reg111 <= $signed((^(&(+((8'haa) != reg97)))));
    end
  assign wire112 = (|reg98[(4'hb):(3'h7)]);
  assign wire113 = $signed(wire70);
  assign wire114 = (+reg80[(4'hd):(1'h1)]);
  assign wire115 = $signed(reg101);
  always
    @(posedge clk) begin
      reg116 <= ({$unsigned({$unsigned(wire89)})} >> $unsigned(wire112));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module7
#( parameter param40 = ((~^{(((8'hb7) < (8'hac)) ~^ (&(8'haf)))}) == ({(~|{(8'ha8), (8'h9d)})} ? {((~|(7'h43)) ? ((8'hb5) ? (8'ha7) : (8'ha6)) : ((8'h9e) & (8'had)))} : ((((8'h9e) ? (7'h40) : (7'h43)) * {(8'had)}) ? (((8'hbe) ? (8'hb7) : (8'ha3)) + ((8'h9d) & (8'hb0))) : {((8'hb3) && (8'hb7)), {(8'hb9), (8'h9e)}}))) )
(y, clk, wire8, wire9, wire10, wire11, wire12);
  output wire [(32'hd2):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h7):(1'h0)] wire8;
  input wire signed [(4'he):(1'h0)] wire9;
  input wire [(4'he):(1'h0)] wire10;
  input wire signed [(5'h15):(1'h0)] wire11;
  input wire signed [(5'h12):(1'h0)] wire12;
  wire signed [(4'h8):(1'h0)] wire39;
  wire [(4'hf):(1'h0)] wire13;
  wire [(5'h14):(1'h0)] wire14;
  wire [(3'h6):(1'h0)] wire15;
  wire [(5'h14):(1'h0)] wire16;
  wire signed [(5'h10):(1'h0)] wire17;
  reg signed [(2'h3):(1'h0)] reg18 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire19;
  wire signed [(5'h14):(1'h0)] wire20;
  wire [(4'h9):(1'h0)] wire21;
  wire [(4'hc):(1'h0)] wire22;
  wire [(5'h15):(1'h0)] wire23;
  wire [(5'h15):(1'h0)] wire24;
  wire signed [(4'hf):(1'h0)] wire25;
  wire [(4'hc):(1'h0)] wire37;
  assign y = {wire39,
                 wire13,
                 wire14,
                 wire15,
                 wire16,
                 wire17,
                 reg18,
                 wire19,
                 wire20,
                 wire21,
                 wire22,
                 wire23,
                 wire24,
                 wire25,
                 wire37,
                 (1'h0)};
  assign wire13 = ($unsigned(({wire11,
                          (^~(8'hbd))} & ((wire11 >> wire12) == (wire9 ?
                          wire12 : (8'hb1))))) ?
                      ({((wire12 ? wire9 : wire12) ?
                              $signed((8'hb0)) : (wire12 < (8'hbc))),
                          (wire12[(3'h6):(1'h0)] | (wire8 <<< (7'h40)))} + $unsigned(((!wire11) ?
                          (wire8 && wire12) : wire9))) : (|wire10[(3'h7):(3'h7)]));
  assign wire14 = $unsigned(($unsigned((8'hb1)) | wire12[(5'h12):(2'h3)]));
  assign wire15 = wire8;
  assign wire16 = (-({wire13} ?
                      $unsigned($unsigned(wire8)) : $unsigned($signed(wire9))));
  assign wire17 = (~|wire10[(4'h8):(3'h5)]);
  always
    @(posedge clk) begin
      reg18 <= wire8[(1'h1):(1'h1)];
    end
  assign wire19 = wire10;
  assign wire20 = (^~(wire17[(4'hd):(1'h1)] ?
                      (wire19 ? wire15 : wire13) : $signed({(-wire16)})));
  assign wire21 = wire20[(5'h14):(3'h6)];
  assign wire22 = wire11;
  assign wire23 = (8'hbb);
  assign wire24 = wire14[(4'h8):(3'h5)];
  assign wire25 = wire11;
  module26 modinst38 (.wire27(wire17), .y(wire37), .clk(clk), .wire28(wire24), .wire29(wire16), .wire31(wire14), .wire30(wire13));
  assign wire39 = (-$signed(wire19[(4'h9):(4'h9)]));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module26  (y, clk, wire31, wire30, wire29, wire28, wire27);
  output wire [(32'h32):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire31;
  input wire [(4'hf):(1'h0)] wire30;
  input wire signed [(2'h3):(1'h0)] wire29;
  input wire signed [(5'h15):(1'h0)] wire28;
  input wire signed [(2'h3):(1'h0)] wire27;
  wire signed [(4'h9):(1'h0)] wire36;
  wire signed [(4'hb):(1'h0)] wire35;
  wire [(2'h3):(1'h0)] wire34;
  wire [(5'h11):(1'h0)] wire33;
  wire signed [(4'h9):(1'h0)] wire32;
  assign y = {wire36, wire35, wire34, wire33, wire32, (1'h0)};
  assign wire32 = $unsigned((8'hb3));
  assign wire33 = {wire27[(2'h3):(1'h0)]};
  assign wire34 = (8'ha8);
  assign wire35 = ($unsigned($signed(($signed(wire27) ?
                          wire29 : ((8'haf) ? wire34 : wire34)))) ?
                      (wire32[(4'h9):(4'h9)] ^ ((-$unsigned(wire32)) ?
                          ((~wire29) <= {wire30,
                              wire33}) : ($unsigned(wire31) || (~&(8'ha6))))) : wire28[(3'h5):(3'h5)]);
  assign wire36 = wire30[(4'h9):(1'h0)];
endmodule