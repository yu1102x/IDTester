module top  (y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'hbf):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h12):(1'h0)] wire0;
  input wire signed [(4'hf):(1'h0)] wire1;
  input wire signed [(5'h13):(1'h0)] wire2;
  input wire signed [(5'h14):(1'h0)] wire3;
  input wire [(4'h8):(1'h0)] wire4;
  wire signed [(4'h9):(1'h0)] wire305;
  wire signed [(3'h5):(1'h0)] wire304;
  wire signed [(4'ha):(1'h0)] wire303;
  wire signed [(5'h15):(1'h0)] wire301;
  reg signed [(5'h11):(1'h0)] reg165 = (1'h0);
  reg [(4'h9):(1'h0)] reg164 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg163 = (1'h0);
  reg [(5'h13):(1'h0)] reg162 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg161 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg160 = (1'h0);
  reg [(4'h8):(1'h0)] reg159 = (1'h0);
  reg [(4'hb):(1'h0)] reg158 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire5;
  wire [(5'h10):(1'h0)] wire6;
  wire signed [(4'hf):(1'h0)] wire156;
  assign y = {wire305,
                 wire304,
                 wire303,
                 wire301,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 wire5,
                 wire6,
                 wire156,
                 (1'h0)};
  assign wire5 = wire3;
  assign wire6 = $unsigned((wire0 ?
                     wire2[(4'hc):(1'h0)] : $signed($unsigned($signed(wire1)))));
  module7 modinst157 (.wire9(wire5), .wire8(wire3), .y(wire156), .wire12(wire2), .wire11(wire1), .clk(clk), .wire10(wire0));
  always
    @(posedge clk) begin
      if ((^($unsigned((|(~wire156))) && {(8'haf)})))
        begin
          reg158 <= $unsigned($unsigned((8'hb7)));
          if (wire4[(1'h0):(1'h0)])
            begin
              reg159 <= $unsigned({$signed($signed((wire4 ? wire4 : wire2)))});
              reg160 <= $signed(wire156);
              reg161 <= ((^~wire2[(3'h4):(2'h2)]) | $unsigned(({$unsigned(wire0)} - ((wire156 ?
                  wire6 : wire3) <<< wire5))));
              reg162 <= ($signed((~$signed((wire5 && wire6)))) ?
                  wire6 : wire0[(4'h9):(3'h4)]);
            end
          else
            begin
              reg159 <= $unsigned($signed((&(8'h9c))));
              reg160 <= $signed(wire0[(3'h7):(3'h4)]);
              reg161 <= $unsigned($signed({(^$signed(reg161)),
                  wire3[(4'hd):(4'ha)]}));
            end
          reg163 <= {{($unsigned((wire0 * reg158)) ?
                      wire6[(4'h8):(2'h3)] : ((~|wire156) ?
                          {(8'ha9)} : wire1[(2'h2):(1'h0)])),
                  {(~&(~|wire6))}}};
          reg164 <= wire6;
        end
      else
        begin
          reg158 <= ($unsigned($signed(reg164)) ?
              wire156 : $signed((~|$unsigned($unsigned((8'hb6))))));
          reg159 <= $signed(wire1[(4'he):(4'h9)]);
        end
      reg165 <= {(reg158 ^~ (((reg162 ^~ (8'ha2)) ?
              (wire156 != wire3) : wire156) | (reg162[(3'h6):(3'h5)] + reg164)))};
    end
  module166 modinst302 (wire301, clk, reg158, reg165, wire156, reg161);
  assign wire303 = $unsigned(wire5);
  assign wire304 = (wire6 ? wire0[(3'h6):(1'h0)] : reg163[(3'h4):(1'h0)]);
  assign wire305 = ($unsigned($unsigned($unsigned(reg163))) | ($signed((~&wire3[(3'h5):(3'h5)])) ^~ $unsigned((8'hb3))));
endmodule

module module166  (y, clk, wire170, wire169, wire168, wire167);
  output wire [(32'h39e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire170;
  input wire [(5'h11):(1'h0)] wire169;
  input wire [(4'hf):(1'h0)] wire168;
  input wire signed [(3'h5):(1'h0)] wire167;
  wire signed [(5'h10):(1'h0)] wire300;
  wire [(2'h2):(1'h0)] wire299;
  reg [(2'h3):(1'h0)] reg298 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg297 = (1'h0);
  reg [(2'h2):(1'h0)] reg296 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg295 = (1'h0);
  reg [(2'h3):(1'h0)] reg294 = (1'h0);
  reg [(5'h13):(1'h0)] reg293 = (1'h0);
  reg [(4'hb):(1'h0)] reg292 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg291 = (1'h0);
  reg [(5'h15):(1'h0)] reg290 = (1'h0);
  reg [(4'ha):(1'h0)] reg289 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg288 = (1'h0);
  reg [(3'h6):(1'h0)] reg287 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg286 = (1'h0);
  reg [(4'h9):(1'h0)] reg285 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg284 = (1'h0);
  reg [(4'hd):(1'h0)] reg283 = (1'h0);
  reg [(5'h10):(1'h0)] reg282 = (1'h0);
  reg [(3'h6):(1'h0)] reg281 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire238;
  reg [(3'h5):(1'h0)] reg216 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg215 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg214 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg213 = (1'h0);
  reg [(2'h3):(1'h0)] reg212 = (1'h0);
  reg [(5'h11):(1'h0)] reg211 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg210 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg209 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg208 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg207 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg206 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg205 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg204 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg203 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire202;
  wire [(4'h9):(1'h0)] wire201;
  wire [(4'hf):(1'h0)] wire200;
  wire signed [(5'h11):(1'h0)] wire199;
  reg [(5'h13):(1'h0)] reg198 = (1'h0);
  reg [(5'h12):(1'h0)] reg197 = (1'h0);
  reg [(5'h15):(1'h0)] reg196 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg195 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg194 = (1'h0);
  reg [(3'h7):(1'h0)] reg193 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg192 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg191 = (1'h0);
  reg [(5'h13):(1'h0)] reg190 = (1'h0);
  reg [(5'h15):(1'h0)] reg189 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg188 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg187 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg186 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg185 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg184 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg183 = (1'h0);
  reg [(3'h5):(1'h0)] reg182 = (1'h0);
  reg [(5'h12):(1'h0)] reg181 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg180 = (1'h0);
  reg [(4'hc):(1'h0)] reg179 = (1'h0);
  reg [(5'h12):(1'h0)] reg178 = (1'h0);
  wire [(3'h5):(1'h0)] wire177;
  wire signed [(5'h13):(1'h0)] wire176;
  wire [(5'h15):(1'h0)] wire175;
  wire [(4'he):(1'h0)] wire174;
  wire [(4'hd):(1'h0)] wire173;
  wire signed [(5'h13):(1'h0)] wire172;
  wire signed [(5'h10):(1'h0)] wire171;
  wire signed [(3'h7):(1'h0)] wire240;
  wire [(3'h4):(1'h0)] wire241;
  wire signed [(3'h7):(1'h0)] wire242;
  wire [(5'h14):(1'h0)] wire279;
  assign y = {wire300,
                 wire299,
                 reg298,
                 reg297,
                 reg296,
                 reg295,
                 reg294,
                 reg293,
                 reg292,
                 reg291,
                 reg290,
                 reg289,
                 reg288,
                 reg287,
                 reg286,
                 reg285,
                 reg284,
                 reg283,
                 reg282,
                 reg281,
                 wire238,
                 reg216,
                 reg215,
                 reg214,
                 reg213,
                 reg212,
                 reg211,
                 reg210,
                 reg209,
                 reg208,
                 reg207,
                 reg206,
                 reg205,
                 reg204,
                 reg203,
                 wire202,
                 wire201,
                 wire200,
                 wire199,
                 reg198,
                 reg197,
                 reg196,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 reg191,
                 reg190,
                 reg189,
                 reg188,
                 reg187,
                 reg186,
                 reg185,
                 reg184,
                 reg183,
                 reg182,
                 reg181,
                 reg180,
                 reg179,
                 reg178,
                 wire177,
                 wire176,
                 wire175,
                 wire174,
                 wire173,
                 wire172,
                 wire171,
                 wire240,
                 wire241,
                 wire242,
                 wire279,
                 (1'h0)};
  assign wire171 = $unsigned($signed($unsigned(((wire169 ^ wire167) & (~&wire168)))));
  assign wire172 = wire170;
  assign wire173 = wire171[(2'h2):(1'h1)];
  assign wire174 = $signed((|$unsigned(($unsigned(wire173) ?
                       $unsigned(wire169) : $unsigned(wire173)))));
  assign wire175 = (((!(~^wire169)) * ((~^(wire172 ? wire173 : wire170)) ?
                       ((wire170 ? wire169 : (8'ha0)) ?
                           wire172[(4'he):(3'h7)] : {wire173,
                               (8'hbf)}) : wire168)) >> ($unsigned(wire169) ?
                       (~|($unsigned((8'ha5)) ?
                           ((8'hb5) ~^ wire168) : (wire167 ?
                               (8'hac) : wire174))) : $signed(((wire172 ?
                           wire168 : wire172) < (wire169 || wire167)))));
  assign wire176 = (+wire169[(4'hf):(2'h2)]);
  assign wire177 = ((~$unsigned({{(8'hb3)}, $unsigned(wire174)})) ?
                       (~wire168[(1'h0):(1'h0)]) : wire173);
  always
    @(posedge clk) begin
      reg178 <= $signed((wire174 ?
          wire174[(4'hb):(4'h8)] : {(&$signed(wire171)),
              (+(wire170 ~^ wire169))}));
      if (($signed($unsigned(((wire173 | wire172) == wire170))) ?
          $signed(($signed($signed((8'hbd))) - ($signed(wire171) ?
              {wire170} : wire173[(2'h3):(1'h0)]))) : $signed(wire172[(1'h1):(1'h1)])))
        begin
          reg179 <= wire171;
          if ((8'hb1))
            begin
              reg180 <= ((~((|wire171[(5'h10):(4'hf)]) >= wire167)) * $signed($signed((reg179 | (^~wire175)))));
              reg181 <= (wire168 ?
                  ($signed(wire167[(3'h5):(3'h5)]) ?
                      wire171 : ({(+reg179), (8'ha6)} ?
                          (^(wire176 < wire176)) : $unsigned(reg179[(3'h7):(1'h0)]))) : ((^wire167[(1'h1):(1'h0)]) ?
                      (^$signed({wire171})) : (($unsigned(wire169) ?
                              reg178[(4'hc):(3'h5)] : $unsigned(wire168)) ?
                          ((reg178 ^ reg180) <= wire174[(3'h4):(1'h0)]) : ($unsigned(reg178) << reg178))));
              reg182 <= wire173;
              reg183 <= $unsigned((wire171 ? $unsigned(reg180) : wire177));
              reg184 <= wire172;
            end
          else
            begin
              reg180 <= $signed((~$unsigned(((wire167 & wire177) && wire176))));
              reg181 <= ((^~(reg178[(5'h10):(4'hc)] ?
                  reg181 : (!(!reg180)))) < (~&(8'ha8)));
              reg182 <= wire175;
            end
          reg185 <= (~(reg184[(4'hb):(2'h3)] - (~wire173[(4'h8):(3'h5)])));
        end
      else
        begin
          reg179 <= wire170[(3'h7):(3'h4)];
          if ((+$signed(wire167[(3'h5):(2'h2)])))
            begin
              reg180 <= $signed($signed($signed((~$signed((8'h9c))))));
              reg181 <= ((((|(~|reg180)) ?
                      (wire176 ?
                          (wire167 <<< reg185) : (!(7'h40))) : {reg178[(4'h9):(4'h9)]}) & reg183) ?
                  (~^(^~($unsigned(reg185) - $unsigned(reg183)))) : reg182);
              reg182 <= $unsigned(((((wire174 + reg184) ?
                      reg181 : $signed(reg180)) ?
                  wire174 : wire172[(3'h5):(3'h5)]) > (wire174[(3'h7):(2'h2)] ^ ($unsigned(reg185) ?
                  (reg182 ~^ wire173) : $unsigned(reg183)))));
              reg183 <= (^(($unsigned((wire172 == reg178)) >>> {{reg184},
                  $signed(wire175)}) && (wire169[(5'h10):(3'h4)] >= wire171)));
            end
          else
            begin
              reg180 <= reg178;
              reg181 <= $unsigned((~^reg178[(5'h12):(4'hc)]));
              reg182 <= wire168;
              reg183 <= (&(wire175[(4'hd):(2'h3)] ?
                  $signed($unsigned((wire174 || reg184))) : wire174));
            end
          reg184 <= reg182[(2'h3):(2'h3)];
        end
      reg186 <= (reg181[(1'h1):(1'h1)] >= reg180);
      reg187 <= {(+(wire173[(4'ha):(3'h4)] ?
              $signed($signed(wire171)) : ((&reg185) ?
                  reg186[(4'hc):(1'h1)] : $unsigned(wire175)))),
          {$signed(((wire177 < (8'hb6)) ^ reg184[(1'h0):(1'h0)])),
              $signed($unsigned($unsigned(wire174)))}};
      if (reg179[(2'h2):(1'h0)])
        begin
          reg188 <= reg184[(4'h8):(2'h2)];
          if ((|reg181))
            begin
              reg189 <= (reg182 ?
                  $unsigned({((wire177 ? (8'h9e) : reg188) ?
                          (wire174 ?
                              wire168 : wire168) : wire167)}) : $unsigned($signed((~&wire177[(3'h4):(2'h2)]))));
              reg190 <= $unsigned(((8'hbc) ?
                  (({reg179, wire172} ? $unsigned(wire171) : wire177) ?
                      wire167[(3'h4):(1'h0)] : ((~wire169) || (+wire174))) : (+$unsigned($unsigned(reg189)))));
              reg191 <= ((|(((reg188 ?
                      reg190 : (8'h9d)) * (reg190 >> reg185)) <= reg190)) ?
                  ((~&reg186[(4'he):(3'h7)]) + $signed($signed(reg188))) : reg184[(2'h2):(1'h1)]);
            end
          else
            begin
              reg189 <= $unsigned(((({reg188} ?
                      (|reg180) : $unsigned(wire169)) ^ $unsigned({reg188})) ?
                  $unsigned($unsigned((reg182 | reg191))) : wire174[(2'h2):(1'h1)]));
              reg190 <= wire175;
              reg191 <= wire172;
              reg192 <= (&$unsigned(wire171[(4'h8):(2'h3)]));
            end
          reg193 <= (|(^(wire173 <<< {reg186[(5'h11):(2'h3)],
              (wire172 ? reg192 : wire177)})));
          reg194 <= reg193;
          if ((8'hba))
            begin
              reg195 <= $signed((^~{(~^$unsigned(reg184)), wire173}));
              reg196 <= wire169;
              reg197 <= ((+reg190[(5'h10):(4'h8)]) ?
                  $unsigned(wire171[(3'h5):(3'h4)]) : $signed((!reg196)));
            end
          else
            begin
              reg195 <= {$signed($unsigned((~|reg193))),
                  (reg179[(4'h8):(2'h2)] ~^ (reg180[(1'h1):(1'h0)] ?
                      ((~(8'hb5)) > reg182) : (reg197[(1'h1):(1'h0)] ?
                          (wire171 ? reg185 : reg192) : {reg186})))};
              reg196 <= $unsigned($unsigned($unsigned((^(~|reg178)))));
              reg197 <= {(&{wire176[(5'h11):(1'h0)], reg191[(3'h5):(1'h1)]})};
              reg198 <= (|$signed($unsigned($unsigned((~|wire167)))));
            end
        end
      else
        begin
          reg188 <= reg195[(2'h2):(1'h1)];
          reg189 <= ($unsigned(reg196[(4'hc):(4'hb)]) ?
              wire171[(4'ha):(2'h2)] : {($signed((reg192 == wire177)) >= wire170),
                  $unsigned($unsigned((wire176 <<< reg189)))});
          if (((reg180[(5'h12):(5'h12)] ?
                  ((reg188[(4'h8):(2'h2)] > reg181) ?
                      ($unsigned((8'ha5)) <<< wire172) : $signed($unsigned(reg183))) : (~^($unsigned(wire167) ?
                      $signed(reg179) : $unsigned(reg179)))) ?
              reg196[(4'he):(4'h8)] : $signed((wire171[(1'h0):(1'h0)] ?
                  reg195[(2'h2):(1'h0)] : wire175[(4'ha):(4'ha)]))))
            begin
              reg190 <= wire167;
              reg191 <= wire175;
            end
          else
            begin
              reg190 <= ($unsigned((reg198 < ($signed(wire176) - (wire168 ?
                  reg185 : reg184)))) == $unsigned((^((^~reg181) ?
                  (8'ha3) : wire172[(5'h11):(4'hd)]))));
              reg191 <= $unsigned($unsigned(reg193[(2'h3):(1'h0)]));
              reg192 <= ({($unsigned((~&wire171)) ?
                      $signed((~(8'ha6))) : (reg185 ? wire172 : (+(8'ha0)))),
                  (8'hb7)} * $unsigned($unsigned($signed((wire170 ?
                  reg178 : reg192)))));
              reg193 <= $unsigned((~|$signed($unsigned((8'hb2)))));
              reg194 <= (reg187[(4'hd):(1'h0)] ?
                  $signed((!reg188[(3'h6):(3'h6)])) : $unsigned(reg192));
            end
          reg195 <= (reg187[(4'hb):(3'h5)] << $signed((wire171[(4'h8):(2'h3)] <<< $signed(reg198))));
          reg196 <= reg197;
        end
    end
  assign wire199 = ((((reg194[(4'he):(3'h4)] ?
                           $unsigned(reg196) : $signed((8'h9e))) ?
                       ($signed(wire177) ?
                           {reg188} : {reg192}) : wire175[(4'hf):(2'h2)]) <= $unsigned(wire173[(1'h1):(1'h1)])) && ((((reg183 ?
                               wire167 : wire177) ?
                           (~^reg187) : (reg182 ^~ reg178)) ?
                       ((reg189 ?
                           reg180 : reg193) ~^ (wire175 >> reg197)) : reg190) <<< {((reg182 > wire170) ?
                           $signed(wire169) : (reg187 >> wire173))}));
  assign wire200 = wire167;
  assign wire201 = ((~|$unsigned($unsigned($signed(reg188)))) ?
                       reg197 : $signed(((reg192[(4'h8):(3'h7)] ?
                               $unsigned(wire168) : (reg198 ?
                                   (8'ha7) : reg178)) ?
                           {(|reg184)} : $unsigned((reg194 ?
                               (8'ha4) : reg189)))));
  assign wire202 = $signed((^$unsigned(reg197)));
  always
    @(posedge clk) begin
      reg203 <= ($signed($signed((+(^reg184)))) | wire176);
      reg204 <= (((~&(&reg187[(1'h0):(1'h0)])) && reg181[(4'h9):(4'h8)]) ?
          ((!((+(7'h40)) ? reg179 : $signed(wire170))) ?
              (8'hb3) : ((!$signed(wire168)) ?
                  wire176[(1'h0):(1'h0)] : ({reg203} ~^ (reg198 ?
                      reg187 : reg178)))) : (~(~|$unsigned($unsigned(wire200)))));
      reg205 <= (reg186[(3'h4):(2'h2)] << wire177);
      if ($unsigned($signed(reg193[(2'h3):(1'h1)])))
        begin
          reg206 <= (^reg194);
        end
      else
        begin
          if (reg190)
            begin
              reg206 <= (+(({$signed(reg187), (reg195 + wire202)} ?
                      $unsigned(wire167[(1'h0):(1'h0)]) : reg190) ?
                  reg189[(4'he):(3'h4)] : (|(~$signed(wire175)))));
              reg207 <= $signed(wire175);
              reg208 <= (~|reg207);
            end
          else
            begin
              reg206 <= {($signed((((8'hbc) ? reg207 : wire168) ?
                      {reg194} : (~&reg184))) ^~ reg181[(4'ha):(3'h6)]),
                  {$signed($signed((reg194 << wire200))),
                      reg195[(1'h1):(1'h1)]}};
            end
          if (wire169)
            begin
              reg209 <= wire199[(3'h6):(2'h3)];
            end
          else
            begin
              reg209 <= (reg208 ?
                  $signed(reg193[(3'h5):(3'h5)]) : $signed($signed((~(^reg198)))));
            end
          if ((8'hbd))
            begin
              reg210 <= wire169[(3'h6):(1'h0)];
            end
          else
            begin
              reg210 <= ((reg180 << $unsigned((~^(-wire199)))) ?
                  {$unsigned((+(8'hbb))), reg209} : $unsigned((!reg193)));
              reg211 <= $signed(wire168[(3'h4):(3'h4)]);
              reg212 <= reg178;
              reg213 <= ({reg184, $signed({(reg210 != reg185), (~(8'hb7))})} ?
                  ($unsigned(wire170) || reg186) : wire168[(4'hb):(4'ha)]);
              reg214 <= (|$unsigned((^reg179)));
            end
          reg215 <= ($unsigned(((wire174[(4'ha):(2'h3)] ^~ (~reg186)) - reg190)) ?
              wire176[(1'h0):(1'h0)] : ({(~^wire174[(4'h8):(3'h4)])} == (!(((8'ha3) >= (8'ha4)) && $unsigned(reg184)))));
        end
      reg216 <= reg192[(4'ha):(4'h8)];
    end
  module217 modinst239 (wire238, clk, wire176, reg185, wire170, wire171, reg192);
  assign wire240 = $signed((wire177[(1'h0):(1'h0)] ?
                       (reg187[(4'hf):(4'hd)] <<< reg182[(3'h4):(2'h2)]) : ((-{reg181,
                           reg192}) + reg182)));
  assign wire241 = (wire199[(4'hd):(4'hb)] ?
                       (reg189 ?
                           ($unsigned($unsigned((8'hb2))) ?
                               (~|(wire177 ? (8'ha0) : wire240)) : (((8'hb5) ?
                                   (8'hb4) : reg181) <<< {reg211})) : (7'h41)) : {(~&{$unsigned(reg182),
                               reg178[(1'h1):(1'h1)]}),
                           ((reg204[(3'h4):(2'h2)] ^ (reg212 <<< reg214)) >> reg198[(5'h11):(3'h4)])});
  assign wire242 = wire170[(1'h0):(1'h0)];
  module243 modinst280 (.wire248(reg205), .wire247(reg186), .wire244(reg208), .wire245(wire169), .wire246(reg191), .y(wire279), .clk(clk));
  always
    @(posedge clk) begin
      reg281 <= reg216;
      if ($signed((~|$unsigned(wire169[(3'h6):(3'h5)]))))
        begin
          reg282 <= (~((~((reg213 ? reg178 : reg207) & {(8'hbd),
              wire200})) == ($unsigned({(8'ha9), reg190}) ? wire170 : reg216)));
          if ((((wire167 ? reg195 : (&(reg193 ? reg186 : (8'hb4)))) ?
              (8'ha5) : $signed((8'ha5))) | (8'hae)))
            begin
              reg283 <= $signed($unsigned(reg182));
              reg284 <= (8'ha7);
              reg285 <= (8'hba);
            end
          else
            begin
              reg283 <= (~$signed($signed(wire176[(5'h13):(2'h2)])));
            end
          reg286 <= $signed(wire170);
          reg287 <= wire170[(3'h5):(3'h5)];
          reg288 <= (&(wire238 ?
              reg203[(3'h4):(2'h2)] : ((((8'hb0) ?
                  (8'hb6) : (8'hb0)) || (&reg212)) && (~wire240[(1'h1):(1'h0)]))));
        end
      else
        begin
          reg282 <= reg189;
        end
      reg289 <= $signed($signed(reg185));
      if (reg215)
        begin
          if ({(~|reg197), $unsigned({(~(reg287 ? (8'hb0) : reg186))})})
            begin
              reg290 <= reg284[(4'h9):(3'h6)];
              reg291 <= $signed(wire177[(1'h1):(1'h1)]);
              reg292 <= (({((reg205 > (8'had)) <= $signed(reg216))} ?
                      ($signed(reg205[(3'h4):(1'h0)]) ?
                          reg204 : (8'hb5)) : ({{reg197, reg190}} ?
                          ($unsigned(reg210) ~^ wire174[(4'hc):(2'h3)]) : (reg210[(1'h1):(1'h1)] ?
                              reg209 : {wire238}))) ?
                  (^~$unsigned($signed(wire169[(4'hc):(3'h5)]))) : (($signed((reg209 > wire238)) ?
                      {(reg184 ? wire241 : (8'hb3)),
                          $unsigned(reg281)} : ((reg189 >>> (8'hae)) - {(7'h42)})) <<< ((~|(reg193 ?
                      (8'hb2) : wire171)) == reg211)));
              reg293 <= {reg195[(1'h1):(1'h0)]};
            end
          else
            begin
              reg290 <= (^$signed(reg178[(3'h4):(2'h3)]));
              reg291 <= {reg289[(1'h0):(1'h0)], (+(wire201 >> (~wire167)))};
              reg292 <= {$signed(wire172)};
            end
          reg294 <= (wire240 ?
              (-$signed((~reg292[(1'h1):(1'h1)]))) : {{reg281,
                      $unsigned($unsigned(reg216))},
                  (^{(~|reg183)})});
          reg295 <= reg206;
          reg296 <= ((^~reg213[(2'h2):(2'h2)]) <<< wire202[(3'h7):(2'h3)]);
          reg297 <= $unsigned((^((+$signed(wire199)) ?
              $signed((reg204 ^~ wire200)) : reg285[(3'h4):(3'h4)])));
        end
      else
        begin
          reg290 <= wire172[(4'hc):(3'h7)];
          reg291 <= reg289;
          reg292 <= reg179[(2'h2):(1'h0)];
          reg293 <= (wire202[(4'hf):(4'h8)] ?
              (&(~|wire240)) : ($signed((-(reg181 << reg293))) ?
                  $unsigned($signed((reg290 ?
                      reg196 : reg286))) : $signed(((reg193 ^ wire200) ~^ reg178))));
          reg294 <= {$signed({$signed((&reg190)),
                  ((reg183 ? reg205 : reg212) ?
                      $signed(reg291) : (reg189 || reg213))})};
        end
      reg298 <= (reg209[(1'h1):(1'h0)] + $signed((-$unsigned((wire176 - reg212)))));
    end
  assign wire299 = reg193[(3'h5):(1'h0)];
  assign wire300 = $unsigned($signed($signed(reg287)));
endmodule

module module7  (y, clk, wire8, wire9, wire10, wire11, wire12);
  output wire [(32'h127):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire8;
  input wire signed [(3'h4):(1'h0)] wire9;
  input wire signed [(5'h12):(1'h0)] wire10;
  input wire signed [(3'h6):(1'h0)] wire11;
  input wire [(5'h13):(1'h0)] wire12;
  wire signed [(3'h5):(1'h0)] wire155;
  reg [(3'h7):(1'h0)] reg154 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire153;
  wire signed [(5'h13):(1'h0)] wire151;
  wire [(4'he):(1'h0)] wire128;
  wire [(5'h10):(1'h0)] wire127;
  wire [(4'ha):(1'h0)] wire126;
  reg [(5'h11):(1'h0)] reg125 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg124 = (1'h0);
  reg [(5'h12):(1'h0)] reg123 = (1'h0);
  reg [(3'h5):(1'h0)] reg122 = (1'h0);
  reg [(5'h13):(1'h0)] reg121 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg120 = (1'h0);
  reg signed [(4'he):(1'h0)] reg119 = (1'h0);
  reg [(3'h4):(1'h0)] reg118 = (1'h0);
  reg [(3'h4):(1'h0)] reg117 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire116;
  wire [(3'h4):(1'h0)] wire115;
  wire signed [(4'h8):(1'h0)] wire113;
  wire signed [(4'hd):(1'h0)] wire63;
  wire signed [(4'h8):(1'h0)] wire13;
  wire [(3'h5):(1'h0)] wire14;
  wire signed [(5'h15):(1'h0)] wire15;
  wire signed [(5'h12):(1'h0)] wire16;
  wire [(5'h14):(1'h0)] wire61;
  assign y = {wire155,
                 reg154,
                 wire153,
                 wire151,
                 wire128,
                 wire127,
                 wire126,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 reg117,
                 wire116,
                 wire115,
                 wire113,
                 wire63,
                 wire13,
                 wire14,
                 wire15,
                 wire16,
                 wire61,
                 (1'h0)};
  assign wire13 = {wire10[(2'h3):(2'h2)]};
  assign wire14 = ((!$signed(((8'hbf) ? $signed(wire8) : $unsigned(wire10)))) ?
                      ((~&$unsigned($unsigned(wire13))) & wire13[(2'h3):(2'h2)]) : $signed($unsigned(((wire9 ?
                              wire8 : (8'hbf)) ?
                          (8'hbd) : $signed(wire11)))));
  assign wire15 = $signed($unsigned({$unsigned((7'h41))}));
  assign wire16 = $signed(wire12);
  module17 modinst62 (.clk(clk), .wire22(wire9), .y(wire61), .wire18(wire10), .wire19(wire16), .wire21(wire14), .wire20(wire15));
  assign wire63 = wire13;
  module64 modinst114 (wire113, clk, wire16, wire63, wire14, wire10);
  assign wire115 = wire11[(3'h6):(1'h1)];
  assign wire116 = (($unsigned(wire113) | ($signed($signed(wire8)) ~^ {(wire115 ^~ (8'ha6))})) <= {(+($unsigned(wire115) ~^ wire115[(3'h4):(1'h0)])),
                       (8'ha7)});
  always
    @(posedge clk) begin
      if (($unsigned((~|{(!wire13)})) && (wire10 ?
          $unsigned(wire10[(3'h5):(2'h3)]) : (wire12[(3'h5):(2'h3)] ?
              wire115[(1'h1):(1'h1)] : $signed((wire12 ? wire16 : (8'hb6)))))))
        begin
          reg117 <= (&(~|$signed((8'hb8))));
          if (($unsigned(($signed((wire14 - wire14)) && wire61)) ?
              $unsigned($signed((~^(-wire8)))) : $signed(wire8)))
            begin
              reg118 <= {(^~wire13[(1'h0):(1'h0)]),
                  $signed(($unsigned((^wire11)) || $signed($unsigned(wire116))))};
              reg119 <= wire9;
              reg120 <= wire63;
              reg121 <= ((~((~|$signed(wire61)) ? wire13 : (~|wire9))) ?
                  ((($unsigned(reg120) >>> $unsigned(wire61)) ?
                          $signed((^wire11)) : wire16[(2'h2):(1'h0)]) ?
                      {wire10} : (|(wire116 & (reg120 ?
                          reg118 : wire13)))) : (wire16 ?
                      (!{(wire116 != reg120)}) : ($signed($signed(reg119)) ?
                          (&wire61) : $signed(wire113[(1'h1):(1'h0)]))));
            end
          else
            begin
              reg118 <= (~^(~^((wire8 && wire16) ?
                  $unsigned((!wire13)) : {{(7'h41)}, {wire13}})));
              reg119 <= wire15[(5'h11):(4'h9)];
            end
        end
      else
        begin
          reg117 <= wire8;
          if (wire115[(2'h3):(1'h0)])
            begin
              reg118 <= $signed((7'h40));
              reg119 <= (^~$unsigned((8'haa)));
            end
          else
            begin
              reg118 <= $signed($signed($signed($signed((~|reg118)))));
              reg119 <= wire63[(3'h5):(2'h3)];
              reg120 <= {reg117[(2'h3):(1'h1)]};
            end
          reg121 <= (^~($signed((wire61 ? (~|wire116) : wire10)) ?
              {{(wire9 ? wire14 : wire9)},
                  $unsigned($unsigned(reg118))} : ($unsigned($unsigned((8'ha4))) ?
                  (~|{wire10}) : wire16[(2'h3):(2'h3)])));
        end
      reg122 <= (($unsigned(({reg118} == wire15[(1'h0):(1'h0)])) ?
          wire16[(4'hd):(3'h7)] : wire11) | reg119);
    end
  always
    @(posedge clk) begin
      reg123 <= (($unsigned(wire113) - wire61[(3'h7):(1'h0)]) ?
          $unsigned({$unsigned($signed(wire61))}) : (^~wire115));
      reg124 <= {((~((^~(8'hb3)) ? $signed(wire13) : (^(8'h9c)))) ?
              $signed(((wire12 ?
                  (8'hb3) : (8'ha3)) ^~ $unsigned(wire10))) : $signed($unsigned(wire12[(4'hc):(2'h2)]))),
          wire61[(4'he):(3'h4)]};
      reg125 <= (((8'ha8) ?
          (!(&(^~(8'hbb)))) : wire63) <<< (wire115[(3'h4):(2'h3)] ~^ (!($signed(reg123) ?
          (reg124 >> reg123) : ((8'hbf) ? wire8 : (8'ha7))))));
    end
  assign wire126 = reg124;
  assign wire127 = ((&(&$signed((reg121 == wire9)))) ?
                       ((8'h9f) ?
                           wire11[(2'h3):(2'h3)] : (^~(wire113[(4'h8):(4'h8)] ?
                               wire16[(2'h3):(2'h2)] : wire15[(3'h4):(2'h2)]))) : (!(8'hb6)));
  assign wire128 = (|wire63);
  module129 modinst152 (.wire133(wire126), .wire131(wire128), .y(wire151), .wire132(wire8), .clk(clk), .wire130(wire61));
  assign wire153 = wire128;
  always
    @(posedge clk) begin
      reg154 <= (^$unsigned($unsigned(reg125)));
    end
  assign wire155 = reg123;
endmodule

module module129
#( parameter param149 = (((8'ha3) > (8'ha5)) ? (-((((8'hb6) ? (8'hb2) : (8'hbb)) << (8'hbd)) + (~&(!(8'ha8))))) : (((((8'ha7) != (8'ha5)) | (8'hbc)) - (((8'ha3) <= (8'hbf)) << (+(8'ha4)))) ? (((&(8'hbc)) <= ((8'ha7) - (8'hb0))) | (~|((7'h44) ? (8'hba) : (8'ha6)))) : ((((8'had) ? (8'hba) : (8'hbb)) ? ((8'hba) + (8'ha5)) : {(8'ha3), (8'hbc)}) >>> {((8'hbf) | (8'hbf))})))
, parameter param150 = (&(((~|(param149 ? param149 : param149)) ? param149 : param149) - param149)) )
(y, clk, wire133, wire132, wire131, wire130);
  output wire [(32'ha9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire133;
  input wire signed [(5'h14):(1'h0)] wire132;
  input wire signed [(4'he):(1'h0)] wire131;
  input wire [(4'h9):(1'h0)] wire130;
  wire signed [(5'h11):(1'h0)] wire148;
  wire signed [(4'hb):(1'h0)] wire147;
  wire signed [(5'h13):(1'h0)] wire146;
  reg [(3'h5):(1'h0)] reg145 = (1'h0);
  reg [(2'h2):(1'h0)] reg144 = (1'h0);
  reg [(3'h5):(1'h0)] reg143 = (1'h0);
  wire [(4'hd):(1'h0)] wire142;
  wire [(4'ha):(1'h0)] wire141;
  wire [(4'hc):(1'h0)] wire140;
  wire signed [(3'h4):(1'h0)] wire139;
  wire signed [(4'h9):(1'h0)] wire138;
  wire [(3'h5):(1'h0)] wire137;
  wire signed [(4'he):(1'h0)] wire136;
  wire signed [(5'h15):(1'h0)] wire135;
  wire signed [(5'h15):(1'h0)] wire134;
  assign y = {wire148,
                 wire147,
                 wire146,
                 reg145,
                 reg144,
                 reg143,
                 wire142,
                 wire141,
                 wire140,
                 wire139,
                 wire138,
                 wire137,
                 wire136,
                 wire135,
                 wire134,
                 (1'h0)};
  assign wire134 = (8'hb8);
  assign wire135 = (-($unsigned(wire132) << wire130[(2'h3):(1'h0)]));
  assign wire136 = ({{(+$signed(wire130)),
                           (~&(!wire133))}} ^ {(($signed(wire132) ?
                           {wire132} : (wire134 ?
                               wire131 : wire132)) == ((wire133 ?
                           wire132 : wire130) != {wire133}))});
  assign wire137 = $signed($unsigned({($signed(wire133) ?
                           $unsigned(wire133) : (~|wire132)),
                       $unsigned(wire131)}));
  assign wire138 = wire136[(4'h9):(2'h2)];
  assign wire139 = $unsigned(((wire130[(2'h2):(1'h1)] * $signed(wire130)) ?
                       (|({wire131,
                           wire130} > {wire135})) : wire130[(4'h9):(3'h5)]));
  assign wire140 = (wire134 ?
                       ($signed(((wire134 < wire133) ?
                               (wire131 ?
                                   wire135 : wire137) : $signed(wire135))) ?
                           (wire138 != wire131[(1'h0):(1'h0)]) : (~|(!(wire131 ?
                               (8'hb1) : wire138)))) : {($signed((wire133 >= wire134)) >= ((|wire138) ?
                               (|(7'h41)) : (wire131 ? wire130 : wire130))),
                           {wire132[(1'h1):(1'h1)],
                               $signed($unsigned((8'hbb)))}});
  assign wire141 = wire140[(2'h3):(1'h0)];
  assign wire142 = (((|wire131[(4'h9):(2'h3)]) ?
                           $signed({wire139[(1'h1):(1'h1)]}) : (wire134[(4'hb):(1'h0)] ?
                               $signed(wire138) : (!$unsigned((8'hbb))))) ?
                       (-wire136) : wire130[(4'h8):(4'h8)]);
  always
    @(posedge clk) begin
      reg143 <= wire139;
      reg144 <= ($unsigned(wire135) * ($signed({(wire139 ?
                  wire132 : wire134)}) ?
          wire137 : reg143));
      reg145 <= $unsigned(wire137);
    end
  assign wire146 = wire132;
  assign wire147 = (8'h9c);
  assign wire148 = $signed(wire142[(4'ha):(3'h7)]);
endmodule

module module64
#( parameter param112 = ((({((8'haa) ? (8'ha1) : (8'hb1))} ? (((8'hac) <<< (8'h9c)) ^ (8'h9f)) : (8'hb9)) ? {(+((7'h42) == (8'ha4))), ((~^(8'ha5)) << ((8'hbb) >>> (8'ha4)))} : (&(((8'hb6) ? (8'hac) : (8'hbd)) ? {(8'h9f)} : ((7'h43) < (8'ha3))))) ^ (((^~((8'ha7) ? (8'ha3) : (8'hab))) < (&(^(8'h9c)))) ? (+(((8'h9d) << (8'hae)) + ((8'hbb) ? (8'hb4) : (8'ha6)))) : (((7'h43) ? ((8'hb0) ? (8'ha9) : (8'hb3)) : ((8'had) ? (8'hb2) : (8'ha1))) * {(|(8'h9e)), (8'hac)}))) )
(y, clk, wire68, wire67, wire66, wire65);
  output wire [(32'h21c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h2):(1'h0)] wire68;
  input wire signed [(4'ha):(1'h0)] wire67;
  input wire [(3'h4):(1'h0)] wire66;
  input wire signed [(2'h3):(1'h0)] wire65;
  wire signed [(4'hf):(1'h0)] wire111;
  wire [(4'hd):(1'h0)] wire110;
  wire signed [(4'h8):(1'h0)] wire109;
  wire [(5'h12):(1'h0)] wire108;
  wire signed [(3'h6):(1'h0)] wire107;
  wire [(5'h15):(1'h0)] wire106;
  wire [(3'h4):(1'h0)] wire105;
  reg signed [(5'h13):(1'h0)] reg104 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg103 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg102 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire101;
  wire [(3'h6):(1'h0)] wire100;
  wire [(5'h12):(1'h0)] wire99;
  wire [(4'hc):(1'h0)] wire98;
  wire signed [(3'h4):(1'h0)] wire97;
  wire [(4'hb):(1'h0)] wire96;
  wire [(4'hb):(1'h0)] wire95;
  reg signed [(5'h14):(1'h0)] reg94 = (1'h0);
  reg [(2'h2):(1'h0)] reg93 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg92 = (1'h0);
  reg signed [(4'he):(1'h0)] reg91 = (1'h0);
  reg [(4'hf):(1'h0)] reg90 = (1'h0);
  reg [(3'h5):(1'h0)] reg89 = (1'h0);
  reg [(5'h12):(1'h0)] reg88 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg87 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg86 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg85 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg84 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg83 = (1'h0);
  wire [(4'hc):(1'h0)] wire82;
  wire signed [(4'hb):(1'h0)] wire81;
  wire signed [(4'hf):(1'h0)] wire80;
  reg [(4'hf):(1'h0)] reg79 = (1'h0);
  reg [(5'h11):(1'h0)] reg78 = (1'h0);
  reg [(2'h3):(1'h0)] reg77 = (1'h0);
  reg [(5'h13):(1'h0)] reg76 = (1'h0);
  reg [(5'h10):(1'h0)] reg75 = (1'h0);
  reg [(4'ha):(1'h0)] reg74 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg73 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg72 = (1'h0);
  reg [(5'h13):(1'h0)] reg71 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg70 = (1'h0);
  wire [(5'h14):(1'h0)] wire69;
  assign y = {wire111,
                 wire110,
                 wire109,
                 wire108,
                 wire107,
                 wire106,
                 wire105,
                 reg104,
                 reg103,
                 reg102,
                 wire101,
                 wire100,
                 wire99,
                 wire98,
                 wire97,
                 wire96,
                 wire95,
                 reg94,
                 reg93,
                 reg92,
                 reg91,
                 reg90,
                 reg89,
                 reg88,
                 reg87,
                 reg86,
                 reg85,
                 reg84,
                 reg83,
                 wire82,
                 wire81,
                 wire80,
                 reg79,
                 reg78,
                 reg77,
                 reg76,
                 reg75,
                 reg74,
                 reg73,
                 reg72,
                 reg71,
                 reg70,
                 wire69,
                 (1'h0)};
  assign wire69 = wire68;
  always
    @(posedge clk) begin
      reg70 <= (&wire67[(2'h3):(2'h2)]);
      if (((8'ha5) ^ ($signed($unsigned(wire69)) ^~ (wire65[(2'h2):(1'h1)] ^ ((+wire65) ?
          wire66[(3'h4):(2'h2)] : $signed(wire68))))))
        begin
          if ((^{$signed(((reg70 > wire69) ~^ $signed(wire66))),
              $signed(wire69)}))
            begin
              reg71 <= $signed($signed($signed($signed($unsigned(wire68)))));
              reg72 <= (($signed((~&wire68)) ?
                      (wire68 ?
                          reg70[(2'h2):(2'h2)] : $signed((!wire68))) : $unsigned(((reg71 >= wire66) ?
                          (reg70 && wire65) : (reg70 ? wire69 : (8'hb5))))) ?
                  (wire69[(5'h11):(1'h0)] != $unsigned(wire67)) : $unsigned(wire67));
              reg73 <= (-{$unsigned($unsigned({reg72, wire69})),
                  {$signed($signed((8'hb6))), {$signed(reg72)}}});
              reg74 <= reg73;
            end
          else
            begin
              reg71 <= $unsigned(reg71);
              reg72 <= $unsigned((($unsigned($signed(wire69)) > wire69[(5'h14):(5'h13)]) <<< ((reg71[(5'h11):(4'hb)] ?
                  (wire65 >= reg72) : reg74) + (wire69 >= (reg74 ^~ reg71)))));
              reg73 <= $unsigned(((((wire66 != (8'haa)) ?
                          $unsigned(wire69) : wire67[(2'h2):(1'h0)]) ?
                      reg71 : ($signed(reg74) <<< ((8'had) ? wire67 : reg72))) ?
                  $unsigned((wire68 != $unsigned(wire66))) : wire65[(1'h0):(1'h0)]));
            end
          reg75 <= $unsigned($signed(($signed({wire65,
              wire65}) + $signed($unsigned(reg74)))));
          if ($signed((~^wire68[(1'h0):(1'h0)])))
            begin
              reg76 <= (|wire66[(2'h3):(1'h0)]);
              reg77 <= wire69[(5'h14):(4'hf)];
            end
          else
            begin
              reg76 <= reg70[(4'hf):(3'h5)];
              reg77 <= wire65;
              reg78 <= ($unsigned($signed(((reg71 ?
                      wire65 : reg73) >>> (reg77 & wire69)))) ?
                  (((!(reg72 ? wire69 : wire67)) ?
                      reg72 : reg72) - $unsigned((^(reg73 ?
                      reg73 : wire65)))) : {$unsigned((wire68[(1'h0):(1'h0)] ?
                          wire66[(2'h3):(2'h3)] : reg71))});
            end
        end
      else
        begin
          reg71 <= {((reg70 ? reg73 : (^~(reg77 ^~ reg74))) ?
                  {$signed($signed((8'h9f)))} : ((!$unsigned(reg72)) - (|(!wire68)))),
              ($unsigned(((reg70 ?
                  reg78 : wire68) - $signed(wire68))) - ($signed($signed(reg70)) != reg78))};
          if (($signed(reg78[(3'h6):(1'h1)]) > (($unsigned((reg78 ?
                  wire65 : wire66)) + $signed((~^reg74))) ?
              (&((-reg73) ?
                  (~(8'hae)) : (wire69 <<< (7'h40)))) : $unsigned($unsigned((reg73 ?
                  reg71 : wire65))))))
            begin
              reg72 <= ($unsigned((reg78[(4'hc):(3'h6)] ?
                  ((+wire68) > $signed(wire67)) : (^~(^(8'ha8))))) * (&($unsigned((~&reg71)) <<< $signed($unsigned(reg75)))));
              reg73 <= ((((7'h41) ?
                      ((wire67 ?
                          reg78 : reg71) - $signed(wire65)) : $signed($unsigned(reg78))) >> $signed({$unsigned(reg72)})) ?
                  (~^reg71[(4'hf):(3'h5)]) : (~^($unsigned((reg73 >> reg75)) ~^ (|(reg77 ?
                      wire69 : reg74)))));
              reg74 <= reg78[(2'h3):(2'h3)];
              reg75 <= reg78;
            end
          else
            begin
              reg72 <= (($signed(((reg78 | wire68) ^ $signed(reg76))) ?
                      $unsigned($signed($unsigned(reg78))) : (wire68 & $unsigned(wire65))) ?
                  reg73 : ((~^($signed((8'hb1)) >> (reg72 ? reg70 : reg70))) ?
                      $signed($unsigned($signed(reg70))) : $unsigned((^~$signed(reg72)))));
              reg73 <= wire69[(4'hf):(4'hc)];
              reg74 <= ((~|(((~(8'hb0)) ?
                  (^~(8'hb9)) : $unsigned(reg75)) <= $signed({(8'hab)}))) < ((wire67 == {$unsigned(wire67),
                      $signed(wire67)}) ?
                  wire69[(2'h2):(2'h2)] : $signed(reg75[(4'h8):(3'h6)])));
              reg75 <= {$unsigned(({reg72} ? {$unsigned(reg70)} : reg72))};
            end
          reg76 <= ((|(($unsigned(reg70) ? (wire65 - reg74) : reg76) ?
                  ((reg72 ? (8'ha7) : reg74) && (reg74 <= wire65)) : reg75)) ?
              (-(+reg70)) : ({$unsigned(reg75[(4'hc):(3'h5)])} - reg75[(4'hb):(3'h5)]));
          reg77 <= ($signed(reg78) ?
              (^($signed(reg72[(2'h3):(1'h1)]) ?
                  ({reg74} < (~^reg70)) : (reg71[(1'h1):(1'h1)] + wire68[(1'h1):(1'h0)]))) : (reg76[(4'h9):(2'h3)] <<< $unsigned((~wire69))));
          reg78 <= $unsigned($unsigned((!(reg71[(4'hc):(4'h8)] ?
              (|(7'h44)) : {reg76}))));
        end
      reg79 <= $unsigned((~&reg77));
    end
  assign wire80 = (+(~((8'ha8) ? {{reg70, reg75}} : (^~$unsigned(wire67)))));
  assign wire81 = $signed($signed({{$signed(reg78)},
                      (^(reg75 ? wire69 : wire67))}));
  assign wire82 = {($signed($unsigned(wire81)) != $signed(reg72[(3'h6):(1'h0)])),
                      ({$unsigned((reg71 ? reg74 : wire80)),
                          wire80[(4'h9):(1'h1)]} == wire68)};
  always
    @(posedge clk) begin
      if ($signed(wire80[(3'h5):(3'h5)]))
        begin
          reg83 <= reg71;
          reg84 <= reg79[(2'h3):(1'h0)];
        end
      else
        begin
          reg83 <= ((8'hb4) ?
              {({{reg72, reg84}} >> ((reg72 ? (7'h41) : reg75) ?
                      $unsigned(reg73) : (~^wire82)))} : reg79);
          reg84 <= reg75[(4'hb):(2'h2)];
        end
      reg85 <= $unsigned($unsigned($unsigned((8'hbe))));
      reg86 <= ({$unsigned({$unsigned(reg72)})} >>> ((~&$unsigned((wire65 >= wire67))) ?
          (^~{$signed(reg72), wire66[(1'h1):(1'h0)]}) : {($signed((8'h9d)) ?
                  {(8'haa)} : reg71)}));
    end
  always
    @(posedge clk) begin
      if ($unsigned(reg79))
        begin
          reg87 <= $signed($unsigned($signed((+$unsigned((7'h44))))));
          reg88 <= (^~$unsigned((!reg87[(2'h3):(2'h3)])));
          if ((|($unsigned({reg73}) ?
              {(reg86[(3'h4):(3'h4)] >= $unsigned(wire81)),
                  $unsigned(reg78)} : $signed((8'hb4)))))
            begin
              reg89 <= ({$signed(wire69[(3'h7):(3'h6)]),
                      ((wire68[(1'h0):(1'h0)] ^~ {reg77, reg84}) ?
                          (wire69[(3'h6):(1'h1)] ?
                              $signed(reg72) : (~|wire69)) : ((reg78 << reg73) || reg87))} ?
                  {(!(((8'ha8) ? reg79 : reg74) ?
                          (reg71 ?
                              wire68 : wire81) : reg72))} : reg72[(2'h2):(1'h1)]);
              reg90 <= wire81[(2'h2):(2'h2)];
            end
          else
            begin
              reg89 <= $signed((&($signed(reg89[(2'h2):(2'h2)]) > reg90)));
              reg90 <= wire82;
              reg91 <= {(-(reg78 != (~&wire80[(1'h0):(1'h0)])))};
              reg92 <= reg90;
            end
          reg93 <= $signed(($signed(((&(8'ha3)) <<< reg72[(3'h7):(1'h0)])) ?
              (({reg73} ? $unsigned((7'h42)) : {reg78, (8'ha4)}) ?
                  reg75[(4'hd):(4'h9)] : ((wire80 + (8'ha8)) ?
                      (reg77 == wire66) : (reg83 ?
                          wire65 : reg78))) : (~^(~^wire69))));
        end
      else
        begin
          reg87 <= reg87;
        end
      reg94 <= $unsigned((^wire66[(1'h1):(1'h0)]));
    end
  assign wire95 = $signed($unsigned((~(|{reg87, (8'hbd)}))));
  assign wire96 = reg70;
  assign wire97 = (8'hb9);
  assign wire98 = $unsigned((((~|(reg71 >> reg78)) ?
                      $unsigned($unsigned(wire96)) : wire82[(1'h0):(1'h0)]) < wire96[(3'h7):(2'h3)]));
  assign wire99 = ((|reg73[(1'h0):(1'h0)]) ?
                      (-(&wire80)) : ({reg91[(2'h2):(2'h2)]} ?
                          $unsigned(wire96) : $unsigned((((8'ha2) ?
                              wire96 : (8'ha7)) ^~ (reg93 || wire68)))));
  assign wire100 = {($signed((-{reg92, wire80})) ?
                           reg71[(3'h6):(3'h5)] : (reg71 ?
                               (+wire82[(3'h6):(2'h2)]) : (8'hba)))};
  assign wire101 = (~|$unsigned(((~|(wire99 != wire82)) && ({reg78} ?
                       wire100[(3'h4):(1'h1)] : $signed((7'h44))))));
  always
    @(posedge clk) begin
      reg102 <= reg73[(2'h2):(1'h0)];
      reg103 <= (wire95[(3'h4):(1'h0)] ?
          ($signed(wire95) ?
              {$signed($signed(wire67)),
                  (+(wire97 ? wire96 : wire65))} : $signed(({wire69,
                  wire80} != $signed((8'ha0))))) : reg79[(4'hb):(3'h7)]);
      reg104 <= (+((((wire96 || wire69) ?
                  $signed(reg78) : (reg78 ? (8'ha1) : reg75)) ?
              $unsigned(reg73[(3'h4):(1'h1)]) : wire68) ?
          wire101[(4'h8):(3'h4)] : $signed(((reg74 != wire82) >= ((7'h41) ?
              wire101 : (8'hb2))))));
    end
  assign wire105 = (($signed((((8'hb5) ?
                               wire99 : (8'haf)) & reg89[(3'h5):(2'h2)])) ?
                           (~&$signed((reg102 >>> wire98))) : ($unsigned(reg92[(4'h9):(4'h9)]) ?
                               {$signed(reg75)} : reg84[(3'h5):(2'h3)])) ?
                       (($unsigned($unsigned((8'hbc))) | reg84[(4'hd):(4'hd)]) + (((reg87 - reg86) | ((8'ha4) ~^ reg89)) || (8'hbd))) : (($signed(reg84[(2'h3):(1'h1)]) <= (wire100[(3'h5):(2'h3)] < (wire67 ?
                           reg83 : reg88))) ^~ ($signed(reg77[(2'h2):(2'h2)]) <= $unsigned(wire66))));
  assign wire106 = (((-wire81[(2'h3):(1'h0)]) & {$unsigned({reg70, (8'ha9)}),
                           (8'hb6)}) ?
                       $unsigned($signed(reg76)) : $unsigned((~&{(wire97 ?
                               (8'haa) : wire99)})));
  assign wire107 = $unsigned((^~$signed(reg72)));
  assign wire108 = ((($signed($signed(reg75)) >= $unsigned($unsigned(wire99))) ?
                       reg91 : $unsigned((-(reg78 || wire66)))) | reg88[(5'h10):(5'h10)]);
  assign wire109 = (wire100 + (^($unsigned((reg74 >> wire106)) - $unsigned($signed(wire95)))));
  assign wire110 = $signed((reg102[(3'h7):(2'h2)] ?
                       (|wire106[(4'hd):(4'hc)]) : $signed($unsigned((wire65 & wire81)))));
  assign wire111 = (~^$unsigned($unsigned($unsigned((&reg74)))));
endmodule

module module17
#( parameter param59 = ((((((8'haf) ~^ (8'hbf)) ~^ ((8'hb4) ~^ (8'hbc))) ? {((8'ha7) >> (8'hbc))} : (+((8'ha1) ? (8'hbc) : (8'haa)))) ? ((!(~(8'haf))) >> (((8'ha4) ? (8'ha6) : (8'haf)) ? ((8'hab) ? (8'hb1) : (8'h9f)) : (8'hbf))) : (~^((~^(8'hb0)) << ((8'ha0) ? (8'hb4) : (8'hb4))))) ? (~^(((~|(7'h43)) ? (-(8'hb0)) : ((8'h9d) ? (8'ha1) : (8'ha3))) & (8'haf))) : ((|(((8'hbe) ^ (7'h40)) ? ((8'hbc) >> (7'h40)) : ((8'hba) ? (8'ha4) : (8'hbd)))) > (({(8'hb3)} > ((8'hac) ? (8'hb5) : (8'ha5))) << (|((8'ha1) < (8'ha5))))))
, parameter param60 = {(|(((param59 < param59) > param59) == (+(8'hb2)))), ((-(~|((8'had) ? param59 : param59))) != param59)} )
(y, clk, wire22, wire21, wire20, wire19, wire18);
  output wire [(32'h16f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h4):(1'h0)] wire22;
  input wire [(3'h5):(1'h0)] wire21;
  input wire [(5'h14):(1'h0)] wire20;
  input wire [(4'hf):(1'h0)] wire19;
  input wire [(4'h8):(1'h0)] wire18;
  wire signed [(3'h6):(1'h0)] wire58;
  wire [(2'h3):(1'h0)] wire57;
  wire signed [(2'h3):(1'h0)] wire56;
  wire [(5'h10):(1'h0)] wire55;
  wire signed [(4'h8):(1'h0)] wire54;
  wire [(4'ha):(1'h0)] wire53;
  wire [(4'hc):(1'h0)] wire52;
  wire [(3'h6):(1'h0)] wire51;
  wire signed [(4'hd):(1'h0)] wire50;
  wire [(3'h7):(1'h0)] wire49;
  reg [(5'h12):(1'h0)] reg48 = (1'h0);
  wire [(4'hc):(1'h0)] wire47;
  wire [(3'h5):(1'h0)] wire46;
  wire signed [(4'hd):(1'h0)] wire45;
  wire signed [(4'hb):(1'h0)] wire44;
  wire signed [(5'h10):(1'h0)] wire43;
  wire signed [(2'h3):(1'h0)] wire42;
  wire [(2'h3):(1'h0)] wire41;
  wire [(4'hf):(1'h0)] wire40;
  wire [(2'h3):(1'h0)] wire39;
  reg signed [(4'hb):(1'h0)] reg38 = (1'h0);
  reg [(3'h4):(1'h0)] reg37 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg36 = (1'h0);
  reg [(4'hf):(1'h0)] reg35 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg34 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg33 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg32 = (1'h0);
  reg [(3'h7):(1'h0)] reg31 = (1'h0);
  reg [(4'hf):(1'h0)] reg30 = (1'h0);
  reg [(5'h14):(1'h0)] reg29 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg28 = (1'h0);
  reg [(4'h8):(1'h0)] reg27 = (1'h0);
  reg [(3'h7):(1'h0)] reg26 = (1'h0);
  reg [(5'h15):(1'h0)] reg25 = (1'h0);
  reg [(5'h15):(1'h0)] reg24 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire23;
  assign y = {wire58,
                 wire57,
                 wire56,
                 wire55,
                 wire54,
                 wire53,
                 wire52,
                 wire51,
                 wire50,
                 wire49,
                 reg48,
                 wire47,
                 wire46,
                 wire45,
                 wire44,
                 wire43,
                 wire42,
                 wire41,
                 wire40,
                 wire39,
                 reg38,
                 reg37,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 reg32,
                 reg31,
                 reg30,
                 reg29,
                 reg28,
                 reg27,
                 reg26,
                 reg25,
                 reg24,
                 wire23,
                 (1'h0)};
  assign wire23 = (+(&$signed($unsigned($signed((7'h41))))));
  always
    @(posedge clk) begin
      reg24 <= (wire20[(4'ha):(3'h5)] ~^ wire18[(1'h1):(1'h0)]);
      reg25 <= {$unsigned($unsigned($unsigned((reg24 ? wire19 : (7'h44)))))};
      reg26 <= (8'hb2);
      if ((8'hbc))
        begin
          reg27 <= (wire19 <<< (reg25[(3'h6):(3'h4)] ? wire18 : wire20));
          if ($unsigned(reg26[(3'h7):(3'h6)]))
            begin
              reg28 <= $signed(wire22[(2'h2):(2'h2)]);
              reg29 <= {{(((8'hab) << (wire20 && wire19)) <<< {$unsigned(wire23)})},
                  (($signed($signed(reg25)) - wire19[(4'ha):(4'h8)]) <<< (+(-{wire20})))};
              reg30 <= reg28[(1'h1):(1'h1)];
              reg31 <= wire18;
              reg32 <= {$unsigned($unsigned((~(!reg29)))), (8'hbe)};
            end
          else
            begin
              reg28 <= ((~&($unsigned((reg32 >>> reg24)) ?
                  (7'h44) : ($signed(wire18) ^ (!reg32)))) & wire18);
              reg29 <= $unsigned(wire18);
              reg30 <= reg29[(3'h6):(3'h4)];
              reg31 <= $signed((~^reg29[(2'h2):(1'h1)]));
              reg32 <= $unsigned((&reg27[(3'h7):(1'h0)]));
            end
          reg33 <= ($unsigned((^(~&(wire19 ?
              reg26 : wire21)))) > $unsigned(((reg31[(3'h5):(2'h3)] || wire18) > {$unsigned(reg29)})));
          if (reg32)
            begin
              reg34 <= (~reg26[(1'h0):(1'h0)]);
            end
          else
            begin
              reg34 <= wire21[(1'h0):(1'h0)];
              reg35 <= $unsigned($unsigned($signed($unsigned((|wire23)))));
              reg36 <= $unsigned(((~^$unsigned($signed((8'ha5)))) > $unsigned((^~(8'ha6)))));
              reg37 <= reg27[(2'h3):(2'h3)];
            end
        end
      else
        begin
          reg27 <= ({$unsigned((~|reg34[(4'hb):(3'h5)]))} ?
              ($unsigned(wire22) | reg30) : $unsigned((reg25[(4'h8):(3'h7)] ?
                  reg32 : ((&reg27) ~^ (-reg31)))));
        end
      reg38 <= ((($signed((~reg32)) & $unsigned($signed(reg35))) ?
          ($unsigned((wire23 << wire21)) | ($signed(reg24) ^~ wire20)) : ((reg27 ?
              (~|reg29) : (reg24 ?
                  reg30 : reg33)) || ($unsigned(wire18) || wire21[(3'h4):(2'h3)]))) != reg33);
    end
  assign wire39 = (|reg32[(3'h6):(2'h3)]);
  assign wire40 = $unsigned($signed((~reg34)));
  assign wire41 = (+({$signed(reg35[(4'ha):(2'h2)])} ?
                      ((~|{reg28}) ?
                          {$signed(reg25),
                              (-reg38)} : (~(wire18 << (8'ha5)))) : wire18[(1'h1):(1'h0)]));
  assign wire42 = $signed((wire19[(4'hc):(2'h3)] >= $signed((~^(reg25 < (8'ha4))))));
  assign wire43 = wire39[(2'h2):(1'h1)];
  assign wire44 = wire19;
  assign wire45 = $signed(reg26[(3'h4):(2'h2)]);
  assign wire46 = $signed(wire43);
  assign wire47 = $signed(reg35[(4'he):(4'hd)]);
  always
    @(posedge clk) begin
      reg48 <= (8'hb1);
    end
  assign wire49 = $unsigned($unsigned(reg25));
  assign wire50 = $unsigned((8'ha4));
  assign wire51 = $unsigned((wire19[(2'h3):(1'h0)] ?
                      wire39 : wire41[(2'h3):(2'h2)]));
  assign wire52 = reg36[(3'h6):(3'h4)];
  assign wire53 = $unsigned($unsigned(reg35));
  assign wire54 = $signed($signed($signed($unsigned(reg32))));
  assign wire55 = (wire20[(4'hf):(4'he)] ? (8'had) : wire54);
  assign wire56 = (^$unsigned(wire51[(1'h1):(1'h0)]));
  assign wire57 = $unsigned($signed(reg29[(2'h2):(1'h0)]));
  assign wire58 = (&(wire56[(1'h1):(1'h0)] ?
                      ($signed({wire53, (8'hb3)}) ~^ ((wire23 ?
                          reg36 : wire43) >>> reg28[(3'h5):(2'h2)])) : $unsigned((~|$signed(wire57)))));
endmodule

module module243
#( parameter param278 = {{((((7'h44) ? (7'h40) : (8'hb8)) >= {(8'hb6), (8'haa)}) ? (((8'h9f) ^ (8'ha3)) ? ((7'h42) ^ (7'h44)) : (~&(8'hbd))) : ((+(8'h9e)) ? (^~(8'had)) : ((8'h9d) ? (8'hae) : (8'hb7)))), (~&(|((8'ha0) - (8'hb2))))}} )
(y, clk, wire248, wire247, wire246, wire245, wire244);
  output wire [(32'h145):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire248;
  input wire [(5'h13):(1'h0)] wire247;
  input wire signed [(5'h13):(1'h0)] wire246;
  input wire [(4'hc):(1'h0)] wire245;
  input wire signed [(5'h14):(1'h0)] wire244;
  wire [(5'h10):(1'h0)] wire277;
  wire signed [(4'hc):(1'h0)] wire276;
  reg signed [(3'h7):(1'h0)] reg275 = (1'h0);
  reg [(3'h7):(1'h0)] reg274 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg273 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg272 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg271 = (1'h0);
  wire [(4'hf):(1'h0)] wire270;
  wire signed [(5'h10):(1'h0)] wire269;
  wire [(4'hc):(1'h0)] wire268;
  wire signed [(2'h3):(1'h0)] wire267;
  wire [(4'ha):(1'h0)] wire266;
  wire [(4'he):(1'h0)] wire265;
  wire signed [(4'h9):(1'h0)] wire264;
  reg [(5'h15):(1'h0)] reg263 = (1'h0);
  reg [(4'hc):(1'h0)] reg262 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg261 = (1'h0);
  reg [(5'h15):(1'h0)] reg260 = (1'h0);
  reg [(2'h2):(1'h0)] reg259 = (1'h0);
  reg [(5'h11):(1'h0)] reg258 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire257;
  wire [(2'h3):(1'h0)] wire256;
  reg signed [(4'hf):(1'h0)] reg255 = (1'h0);
  reg signed [(4'he):(1'h0)] reg254 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg253 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg252 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire251;
  wire [(4'he):(1'h0)] wire250;
  wire [(3'h5):(1'h0)] wire249;
  assign y = {wire277,
                 wire276,
                 reg275,
                 reg274,
                 reg273,
                 reg272,
                 reg271,
                 wire270,
                 wire269,
                 wire268,
                 wire267,
                 wire266,
                 wire265,
                 wire264,
                 reg263,
                 reg262,
                 reg261,
                 reg260,
                 reg259,
                 reg258,
                 wire257,
                 wire256,
                 reg255,
                 reg254,
                 reg253,
                 reg252,
                 wire251,
                 wire250,
                 wire249,
                 (1'h0)};
  assign wire249 = wire248[(1'h1):(1'h0)];
  assign wire250 = {wire245[(3'h6):(2'h3)]};
  assign wire251 = wire250;
  always
    @(posedge clk) begin
      reg252 <= ((($signed((&wire249)) && {(|wire247),
              {wire244}}) ^~ (~|(8'haa))) ?
          wire250 : (~^wire244[(5'h13):(4'hc)]));
      reg253 <= wire249[(3'h4):(1'h1)];
      reg254 <= ($signed((~^$signed(wire250))) < $unsigned($unsigned($signed((wire251 ?
          (8'ha4) : wire249)))));
      reg255 <= ($unsigned({({wire250,
              (8'ha0)} || wire245)}) >>> (~&wire247[(4'h8):(1'h0)]));
    end
  assign wire256 = reg253[(3'h6):(3'h5)];
  assign wire257 = $signed($signed({(^~{reg253})}));
  always
    @(posedge clk) begin
      reg258 <= wire246[(2'h2):(2'h2)];
      reg259 <= ((-$signed(wire257)) != (reg255 ?
          {wire248,
              $signed(wire251)} : (($signed(reg253) && $unsigned(reg253)) ?
              $unsigned(((8'hb9) ? reg255 : reg252)) : $unsigned((^reg253)))));
    end
  always
    @(posedge clk) begin
      reg260 <= ($unsigned(wire257[(2'h2):(2'h2)]) ?
          wire246[(4'h9):(3'h5)] : wire247[(5'h12):(5'h10)]);
      reg261 <= (({(~|{(7'h43), reg253}), (!$unsigned(wire245))} ?
          $signed($unsigned((reg260 ?
              (8'h9c) : wire251))) : wire251[(3'h4):(3'h4)]) + ((({wire248} - $unsigned((8'h9e))) ?
          wire244 : ((reg258 ~^ wire248) ~^ wire249)) & (~|(~&$unsigned(reg253)))));
      reg262 <= $signed(((wire248[(3'h6):(1'h1)] ?
          (-(reg261 ?
              reg259 : wire246)) : $signed(wire249[(3'h4):(1'h1)])) > (8'h9c)));
      reg263 <= ($unsigned(wire256[(2'h3):(2'h3)]) ?
          wire246 : ({$signed(wire256), $unsigned(wire247)} ?
              wire250 : $signed(({wire257, wire249} ?
                  wire257[(1'h1):(1'h1)] : (~^(8'hb8))))));
    end
  assign wire264 = reg260;
  assign wire265 = {(~&($unsigned({reg261}) ? wire247 : (~^$signed(reg262))))};
  assign wire266 = $signed($unsigned(((^~(wire257 ? reg260 : reg253)) ?
                       (reg254 ?
                           (^reg253) : (~wire247)) : $unsigned((~&(8'hb0))))));
  assign wire267 = {reg263,
                       (($signed(wire256) + reg253[(2'h3):(1'h0)]) ^ $unsigned((^~wire264)))};
  assign wire268 = ((~^reg253[(1'h1):(1'h0)]) << (8'hb5));
  assign wire269 = (8'h9f);
  assign wire270 = (^(($unsigned($unsigned(wire251)) ?
                           (&$unsigned(reg260)) : wire266[(4'ha):(3'h6)]) ?
                       (8'ha6) : $unsigned((wire257 << (wire256 ?
                           reg253 : reg253)))));
  always
    @(posedge clk) begin
      reg271 <= (~|wire257);
      reg272 <= (reg271 ^~ reg263[(2'h2):(2'h2)]);
      reg273 <= $unsigned((wire256 ?
          $unsigned(wire266) : (({wire248} << $unsigned(wire245)) >> wire256)));
      reg274 <= wire268;
      reg275 <= $unsigned($signed((wire267[(2'h3):(2'h3)] ?
          (wire245[(4'h8):(3'h7)] ?
              (wire268 ?
                  reg252 : (8'ha1)) : wire248) : ($unsigned(wire257) & $signed(reg261)))));
    end
  assign wire276 = {(((-wire246) == $signed(reg255)) ^~ wire244[(3'h4):(2'h2)])};
  assign wire277 = (~|{$unsigned(($unsigned(wire256) || reg252[(4'hd):(4'h8)]))});
endmodule

module module217
#( parameter param236 = (7'h41)
, parameter param237 = (({{param236}} ? param236 : param236) >> (-((!(|param236)) - ({(8'ha8), (8'ha8)} ? (param236 == param236) : param236)))) )
(y, clk, wire222, wire221, wire220, wire219, wire218);
  output wire [(32'hb7):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h13):(1'h0)] wire222;
  input wire signed [(2'h2):(1'h0)] wire221;
  input wire [(4'hb):(1'h0)] wire220;
  input wire [(4'hd):(1'h0)] wire219;
  input wire signed [(3'h4):(1'h0)] wire218;
  wire [(5'h15):(1'h0)] wire235;
  wire signed [(4'h9):(1'h0)] wire234;
  wire [(4'hd):(1'h0)] wire233;
  wire signed [(4'he):(1'h0)] wire232;
  wire signed [(4'hd):(1'h0)] wire231;
  wire signed [(5'h11):(1'h0)] wire230;
  wire [(4'h8):(1'h0)] wire229;
  wire signed [(5'h13):(1'h0)] wire228;
  reg signed [(4'hd):(1'h0)] reg227 = (1'h0);
  reg [(5'h15):(1'h0)] reg226 = (1'h0);
  reg [(2'h3):(1'h0)] reg225 = (1'h0);
  reg [(5'h10):(1'h0)] reg224 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire223;
  assign y = {wire235,
                 wire234,
                 wire233,
                 wire232,
                 wire231,
                 wire230,
                 wire229,
                 wire228,
                 reg227,
                 reg226,
                 reg225,
                 reg224,
                 wire223,
                 (1'h0)};
  assign wire223 = (~|$signed(((-(wire219 ^ wire218)) ?
                       $unsigned($signed(wire222)) : ($unsigned(wire222) * (^wire222)))));
  always
    @(posedge clk) begin
      reg224 <= (wire222[(2'h3):(1'h1)] ?
          $signed(wire219) : (wire222[(3'h6):(1'h1)] != ($signed($unsigned(wire218)) ^ wire222[(4'he):(2'h3)])));
      reg225 <= ($unsigned($signed($unsigned($unsigned(wire223)))) ?
          {$signed(wire223)} : $unsigned({((wire222 ? wire220 : wire219) ?
                  (reg224 ? reg224 : (8'hbc)) : (wire218 | reg224))}));
      reg226 <= (wire219 <<< (((8'hb5) * ((~|reg225) ^ (~wire222))) >>> wire220));
      reg227 <= $unsigned((wire218[(3'h4):(2'h3)] < ((&(^~reg226)) ?
          (^wire221) : reg224[(4'he):(4'h8)])));
    end
  assign wire228 = $unsigned(wire223);
  assign wire229 = (~&$unsigned(wire222));
  assign wire230 = (wire221 ?
                       $signed((&$unsigned((&wire220)))) : $signed(wire229[(1'h1):(1'h0)]));
  assign wire231 = $signed($signed((($unsigned(wire223) ?
                           $signed(wire222) : reg226) ?
                       ($signed(reg226) == reg224[(3'h5):(1'h0)]) : (reg226 ?
                           ((8'ha6) * reg224) : reg225[(2'h2):(2'h2)]))));
  assign wire232 = (wire222[(4'h9):(1'h1)] >>> {{reg227[(1'h0):(1'h0)]}});
  assign wire233 = {wire229[(2'h2):(1'h1)], wire223[(1'h0):(1'h0)]};
  assign wire234 = ((($signed((wire218 ^~ wire218)) ?
                           {(reg225 ?
                                   wire229 : wire223)} : ((wire233 & wire232) ?
                               $unsigned((8'hb7)) : $signed(wire231))) ?
                       ({(8'h9d)} ?
                           $unsigned($signed(wire228)) : wire222) : $unsigned(wire231)) + (8'hba));
  assign wire235 = ($signed({(wire234 ^ (~|wire221))}) ?
                       {($unsigned((wire219 ?
                               (8'had) : reg227)) >> ((wire222 ~^ wire228) <<< $signed((8'ha8))))} : wire222);
endmodule