module top_1
#( parameter param257 = {(((((7'h41) ? (8'h9e) : (8'hb3)) ? (~|(7'h44)) : ((8'h9e) ? (8'ha6) : (8'h9f))) ? ((8'hae) & {(8'h9e)}) : (^~((8'hb5) ? (8'hbd) : (8'ha4)))) ? ((8'hac) << ({(7'h43), (7'h40)} ? ((8'hbe) && (8'hb1)) : (~^(8'hb8)))) : ((((8'hab) ? (8'ha4) : (8'h9d)) ? ((7'h41) ? (8'hab) : (8'hb1)) : (|(8'hb9))) & (^~{(8'hb6)}))), (8'hb3)}
, parameter param258 = {(~^param257), (param257 - (-(8'h9d)))} )
(y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h180):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire3;
  input wire [(5'h15):(1'h0)] wire2;
  input wire [(5'h11):(1'h0)] wire1;
  input wire [(5'h15):(1'h0)] wire0;
  wire [(4'hc):(1'h0)] wire256;
  wire [(5'h10):(1'h0)] wire255;
  wire [(3'h6):(1'h0)] wire254;
  reg [(4'hd):(1'h0)] reg253 = (1'h0);
  reg [(3'h6):(1'h0)] reg252 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg251 = (1'h0);
  reg [(3'h7):(1'h0)] reg250 = (1'h0);
  wire [(4'h8):(1'h0)] wire249;
  wire signed [(4'ha):(1'h0)] wire248;
  wire signed [(3'h7):(1'h0)] wire247;
  wire signed [(3'h5):(1'h0)] wire246;
  wire signed [(5'h15):(1'h0)] wire242;
  reg [(3'h4):(1'h0)] reg106 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg105 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg104 = (1'h0);
  reg signed [(4'he):(1'h0)] reg103 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg102 = (1'h0);
  reg [(5'h10):(1'h0)] reg101 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg100 = (1'h0);
  reg [(3'h5):(1'h0)] reg99 = (1'h0);
  reg [(5'h11):(1'h0)] reg98 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg97 = (1'h0);
  reg [(4'hf):(1'h0)] reg96 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg95 = (1'h0);
  reg [(4'ha):(1'h0)] reg94 = (1'h0);
  reg [(5'h10):(1'h0)] reg93 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg92 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire91;
  wire signed [(4'h8):(1'h0)] wire90;
  wire signed [(5'h11):(1'h0)] wire88;
  wire signed [(4'hf):(1'h0)] wire244;
  assign y = {wire256,
                 wire255,
                 wire254,
                 reg253,
                 reg252,
                 reg251,
                 reg250,
                 wire249,
                 wire248,
                 wire247,
                 wire246,
                 wire242,
                 reg106,
                 reg105,
                 reg104,
                 reg103,
                 reg102,
                 reg101,
                 reg100,
                 reg99,
                 reg98,
                 reg97,
                 reg96,
                 reg95,
                 reg94,
                 reg93,
                 reg92,
                 wire91,
                 wire90,
                 wire88,
                 wire244,
                 (1'h0)};
  module4_1 modinst89 (wire88, clk, wire1, wire3, wire0, wire2);
  assign wire90 = $unsigned($unsigned(wire3[(4'h9):(4'h9)]));
  assign wire91 = ($signed((((wire1 ? wire88 : wire88) > {wire90,
                      wire3}) ~^ ($signed(wire2) ?
                      $signed(wire2) : (wire1 ?
                          wire3 : wire2)))) >>> {$signed(wire2[(4'hf):(3'h4)]),
                      wire88});
  always
    @(posedge clk) begin
      reg92 <= {((8'h9c) - $signed($unsigned(wire0[(1'h1):(1'h1)]))),
          $signed(wire1)};
      reg93 <= (~^(^((^wire0[(4'h8):(1'h1)]) ?
          wire2 : $unsigned($signed(wire90)))));
      reg94 <= wire0;
      if ($unsigned($signed($unsigned(((wire0 ? (8'ha3) : wire90) ?
          $unsigned(reg92) : (^reg92))))))
        begin
          if (($unsigned(reg94) <<< (~^(^wire88))))
            begin
              reg95 <= wire2[(4'hf):(1'h0)];
              reg96 <= (^~(^$unsigned(wire90[(3'h6):(2'h3)])));
              reg97 <= wire3[(5'h10):(4'h9)];
              reg98 <= $unsigned({$signed((|$unsigned(reg96)))});
              reg99 <= reg98;
            end
          else
            begin
              reg95 <= ((wire1[(1'h1):(1'h1)] ?
                      {reg95} : ($signed($unsigned(reg96)) <<< reg92[(4'ha):(1'h0)])) ?
                  reg95 : {(!$signed(wire91[(5'h13):(4'hf)]))});
              reg96 <= $signed(($unsigned((^~reg99[(2'h2):(1'h1)])) > ($unsigned((8'had)) ?
                  $unsigned(((8'h9c) >>> reg92)) : {reg99})));
              reg97 <= $signed((reg99[(1'h0):(1'h0)] >> (8'h9c)));
              reg98 <= reg93;
            end
          reg100 <= $unsigned(((~&(wire3 ?
              wire88 : (|reg97))) - (wire88[(5'h10):(4'hd)] || (~^(!wire1)))));
        end
      else
        begin
          if (((^~$signed(((reg100 ~^ (8'ha6)) ?
              (reg96 | reg95) : wire88))) != $unsigned((!reg99))))
            begin
              reg95 <= {$unsigned((wire88[(4'hf):(3'h7)] ?
                      {(wire0 ? reg100 : reg97)} : ((~&wire90) ?
                          (|reg100) : wire90)))};
              reg96 <= $signed({(reg92[(5'h12):(3'h5)] ?
                      ($unsigned(reg100) ?
                          $signed(reg100) : wire90) : (~((8'hbc) ?
                          reg96 : reg98)))});
              reg97 <= $unsigned(reg99);
              reg98 <= (reg95 - (8'had));
              reg99 <= reg100;
            end
          else
            begin
              reg95 <= ((^~reg95[(3'h5):(2'h3)]) ?
                  reg95[(1'h0):(1'h0)] : (wire3[(1'h0):(1'h0)] << wire90));
            end
          reg100 <= reg93[(3'h5):(1'h1)];
          if ({wire90})
            begin
              reg101 <= wire3;
              reg102 <= wire2[(2'h2):(1'h0)];
              reg103 <= ({$unsigned(reg99[(2'h2):(1'h0)]),
                      $unsigned(((reg93 ? reg99 : wire3) ?
                          wire90 : reg94[(2'h2):(1'h0)]))} ?
                  (!$signed((~reg93))) : reg94[(1'h1):(1'h0)]);
            end
          else
            begin
              reg101 <= (reg103[(3'h7):(2'h2)] ^ wire90[(2'h3):(2'h3)]);
              reg102 <= (7'h44);
              reg103 <= wire0;
              reg104 <= $signed((((8'haf) ?
                  wire3[(5'h12):(4'hd)] : $signed((8'hba))) + $unsigned((reg94 ?
                  $signed(reg99) : (8'hbc)))));
            end
          reg105 <= $unsigned(reg102[(4'h8):(3'h4)]);
        end
      reg106 <= $unsigned({$unsigned(((-reg94) ?
              (8'ha0) : (wire0 ? reg103 : reg100)))});
    end
  module107_1 modinst243 (.clk(clk), .wire110(reg102), .y(wire242), .wire111(reg101), .wire108(reg96), .wire109(reg92), .wire112(reg97));
  module107_1 modinst245 (.wire110(reg104), .wire111(reg105), .clk(clk), .wire108(reg103), .y(wire244), .wire112(reg94), .wire109(reg100));
  assign wire246 = $signed((reg104 ?
                       reg98 : ((8'haa) ?
                           $signed((reg102 ? wire88 : (8'hb5))) : wire2)));
  assign wire247 = $signed((reg100 ? wire1 : reg93));
  assign wire248 = (($unsigned(wire246) ?
                       $signed((!(!reg94))) : (reg106[(2'h3):(2'h3)] ?
                           $signed(reg103[(3'h5):(2'h3)]) : {(+(7'h43)),
                               (~|wire244)})) + (~&wire91[(2'h2):(2'h2)]));
  assign wire249 = ($unsigned(wire88) ?
                       $signed((!(8'hbe))) : reg99[(2'h2):(1'h0)]);
  always
    @(posedge clk) begin
      reg250 <= ($signed(((!reg94) >= $signed(reg95))) ?
          $unsigned(wire246[(1'h0):(1'h0)]) : wire242);
      reg251 <= (!$signed((~reg98)));
      reg252 <= $signed(reg250);
      reg253 <= wire249;
    end
  assign wire254 = (($signed(reg93[(4'h9):(4'h8)]) ^~ reg106[(3'h4):(3'h4)]) > ((^(^{wire242,
                           (8'ha1)})) ?
                       (|$signed($signed(wire249))) : ((reg250[(1'h0):(1'h0)] ?
                           $unsigned(wire1) : {wire3,
                               reg100}) >> $unsigned(reg102))));
  assign wire255 = reg93;
  assign wire256 = (wire91[(3'h4):(3'h4)] ? reg97 : reg251);
endmodule

module module107_1
#( parameter param241 = ((|((!(~|(8'ha3))) ? (&(~|(8'h9f))) : {{(8'hac), (8'hac)}})) ? ((({(7'h44), (8'hbd)} << (+(8'ha4))) ? (((8'hb8) ^ (8'h9f)) - {(8'had)}) : (((8'ha6) && (8'hae)) ? (~|(8'ha4)) : (|(8'haf)))) > (({(8'hae), (8'h9d)} <= ((8'haa) + (8'hb9))) ~^ {((8'hb5) ? (8'hb5) : (8'h9f))})) : (&((((8'ha1) || (8'hb3)) ? (|(8'hb1)) : ((8'hbd) || (8'ha9))) ? ((7'h41) <= ((8'hb7) ? (8'hb6) : (8'hac))) : (8'haf)))) )
(y, clk, wire112, wire111, wire110, wire109, wire108);
  output wire [(32'h1dd):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire112;
  input wire signed [(2'h3):(1'h0)] wire111;
  input wire signed [(5'h13):(1'h0)] wire110;
  input wire signed [(4'ha):(1'h0)] wire109;
  input wire [(4'he):(1'h0)] wire108;
  wire [(4'hb):(1'h0)] wire240;
  wire signed [(2'h2):(1'h0)] wire239;
  wire signed [(2'h3):(1'h0)] wire238;
  wire signed [(5'h11):(1'h0)] wire237;
  reg [(5'h12):(1'h0)] reg236 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg235 = (1'h0);
  reg [(4'hc):(1'h0)] reg234 = (1'h0);
  reg [(4'h8):(1'h0)] reg233 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg232 = (1'h0);
  reg [(4'ha):(1'h0)] reg231 = (1'h0);
  reg [(5'h14):(1'h0)] reg230 = (1'h0);
  wire [(5'h12):(1'h0)] wire229;
  reg [(5'h14):(1'h0)] reg228 = (1'h0);
  reg [(5'h13):(1'h0)] reg227 = (1'h0);
  reg [(4'h8):(1'h0)] reg226 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg225 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg224 = (1'h0);
  reg [(3'h5):(1'h0)] reg223 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg222 = (1'h0);
  reg [(4'hc):(1'h0)] reg221 = (1'h0);
  reg [(2'h2):(1'h0)] reg220 = (1'h0);
  wire [(4'h8):(1'h0)] wire219;
  wire [(4'h8):(1'h0)] wire217;
  wire signed [(5'h13):(1'h0)] wire132;
  wire signed [(5'h10):(1'h0)] wire131;
  reg [(4'hd):(1'h0)] reg130 = (1'h0);
  reg [(3'h4):(1'h0)] reg129 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg128 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg127 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg126 = (1'h0);
  reg [(5'h14):(1'h0)] reg125 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg124 = (1'h0);
  reg [(4'h8):(1'h0)] reg123 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg122 = (1'h0);
  reg [(2'h3):(1'h0)] reg121 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg120 = (1'h0);
  reg signed [(4'he):(1'h0)] reg119 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg118 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg117 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg116 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg115 = (1'h0);
  wire [(4'hd):(1'h0)] wire114;
  wire [(3'h7):(1'h0)] wire113;
  assign y = {wire240,
                 wire239,
                 wire238,
                 wire237,
                 reg236,
                 reg235,
                 reg234,
                 reg233,
                 reg232,
                 reg231,
                 reg230,
                 wire229,
                 reg228,
                 reg227,
                 reg226,
                 reg225,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 wire219,
                 wire217,
                 wire132,
                 wire131,
                 reg130,
                 reg129,
                 reg128,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 reg117,
                 reg116,
                 reg115,
                 wire114,
                 wire113,
                 (1'h0)};
  assign wire113 = ((({wire108[(4'hc):(3'h7)]} ?
                           (((8'ha0) ?
                               wire109 : wire109) ^ (wire112 * wire112)) : wire112[(1'h1):(1'h1)]) & {($signed(wire108) ?
                               (wire108 ?
                                   wire110 : wire112) : wire110[(5'h13):(1'h1)])}) ?
                       wire109 : $signed(((wire110 ?
                               {wire109} : wire111[(1'h1):(1'h0)]) ?
                           ($unsigned(wire109) ?
                               $signed(wire108) : (wire110 ?
                                   wire109 : wire112)) : wire108[(4'he):(4'h8)])));
  assign wire114 = wire110;
  always
    @(posedge clk) begin
      reg115 <= $unsigned({$unsigned((~^$unsigned(wire114)))});
      reg116 <= $unsigned(wire113[(3'h4):(1'h0)]);
      if ($signed($unsigned((wire112[(1'h1):(1'h0)] && ({wire108} != $unsigned(reg116))))))
        begin
          reg117 <= $signed($unsigned($signed({(^wire114),
              wire110[(5'h12):(3'h7)]})));
          reg118 <= {reg117, wire113};
          reg119 <= (((7'h42) >> wire113[(3'h5):(1'h0)]) == wire110);
        end
      else
        begin
          if (wire109[(2'h2):(2'h2)])
            begin
              reg117 <= wire113[(3'h6):(1'h1)];
              reg118 <= ($unsigned(reg119[(4'h8):(3'h7)]) <<< (($signed((8'haa)) ?
                      ((wire111 >= reg115) & (reg115 == (7'h44))) : (wire113[(3'h4):(1'h0)] ?
                          wire113 : {reg116})) ?
                  (wire114 - $signed(wire110)) : {(wire112 <<< (8'h9d))}));
            end
          else
            begin
              reg117 <= wire108[(4'ha):(1'h0)];
              reg118 <= $unsigned($unsigned($signed(((reg117 ?
                  wire114 : wire111) <<< (~|wire113)))));
              reg119 <= reg118[(1'h0):(1'h0)];
              reg120 <= reg116;
              reg121 <= ($unsigned($unsigned((((8'hbb) ?
                      wire112 : wire114) && (wire112 >> reg118)))) ?
                  (wire113 == {(~|(wire112 ?
                          wire112 : reg117))}) : ($signed(reg119[(4'hb):(3'h4)]) >>> $unsigned((wire114[(4'hc):(1'h1)] ?
                      (wire109 ? reg119 : reg116) : $signed((7'h42))))));
            end
          reg122 <= ($signed({wire111, (|reg118)}) >>> (wire109[(1'h1):(1'h1)] ?
              (~^($unsigned(wire108) ?
                  $signed(wire108) : wire109)) : reg121[(2'h2):(1'h0)]));
          reg123 <= ((|$signed(wire111)) | wire112);
          reg124 <= $signed((((~&wire110[(4'h9):(3'h4)]) - ($signed(wire111) ^ $signed(wire109))) ?
              (((reg117 * (7'h40)) & {reg115, reg121}) ?
                  reg123[(2'h3):(1'h1)] : wire111[(2'h3):(1'h1)]) : reg121[(2'h2):(2'h2)]));
          reg125 <= (wire112[(2'h3):(2'h2)] & ({reg121} ?
              $signed({{wire109, reg122}}) : reg119[(4'ha):(2'h3)]));
        end
      if (((+(~|($unsigned(reg121) > wire110[(4'hf):(2'h2)]))) ?
          $unsigned((~^(|(8'h9f)))) : reg125))
        begin
          reg126 <= reg121[(2'h3):(2'h3)];
          if ((wire110 ?
              (($unsigned($unsigned(reg120)) ?
                      (+(reg123 ~^ reg120)) : reg119[(2'h3):(1'h1)]) ?
                  $signed((~&(~&(8'hb2)))) : $signed(reg118)) : ((reg125 - (wire114 | {reg122,
                  reg123})) & {reg118[(3'h6):(2'h3)]})))
            begin
              reg127 <= {$unsigned(($signed(reg120[(3'h7):(3'h5)]) ?
                      reg121 : $unsigned((^~reg124))))};
              reg128 <= $signed(($signed(((wire112 >>> wire113) ?
                      {reg119} : $unsigned(reg124))) ?
                  $signed($signed($signed(wire110))) : (wire108[(4'h8):(1'h1)] | $signed($signed((8'hae))))));
              reg129 <= ((wire110[(2'h2):(1'h1)] >= (wire114[(4'h9):(1'h0)] ?
                  ((reg124 ~^ wire114) ~^ {reg127,
                      wire110}) : {reg117[(5'h10):(4'h8)],
                      (~|wire111)})) ^~ ($unsigned(reg125) == $signed(reg120[(3'h4):(1'h1)])));
              reg130 <= reg128;
            end
          else
            begin
              reg127 <= $signed((reg116[(4'h8):(1'h0)] ?
                  {(&$signed(reg122))} : $signed(wire114)));
              reg128 <= ($unsigned(((reg123 < $unsigned(wire111)) ?
                      ((&(8'had)) ?
                          reg126[(2'h2):(2'h2)] : (wire108 > wire110)) : ((+reg117) - $unsigned(wire110)))) ?
                  (^reg119[(2'h2):(2'h2)]) : (~(^(reg128 - $unsigned(reg116)))));
            end
        end
      else
        begin
          reg126 <= {$unsigned((~$signed($unsigned(reg129)))),
              $signed(((reg121 != wire111[(1'h1):(1'h1)]) ?
                  ($unsigned(wire109) ?
                      {reg125} : ((8'hbd) ? (8'haa) : wire113)) : ((&reg116) ?
                      (wire109 - wire113) : (reg117 ? reg128 : (8'hb1)))))};
        end
    end
  assign wire131 = reg120[(2'h3):(2'h3)];
  assign wire132 = ((!reg119[(1'h0):(1'h0)]) ?
                       (((reg120[(5'h10):(4'hd)] <= {reg125}) ?
                               ($signed(wire109) ?
                                   reg130 : reg119[(4'hd):(3'h6)]) : {((8'ha0) || reg127),
                                   $signed((8'hb7))}) ?
                           (&$unsigned(reg116[(4'hb):(3'h7)])) : $signed($signed((wire109 & (7'h43))))) : $unsigned($signed(reg117)));
  module133_1 modinst218 (wire217, clk, wire108, reg126, reg118, reg130);
  assign wire219 = (~{wire217[(4'h8):(3'h7)],
                       $signed(((~|(8'hba)) != (reg115 && (7'h43))))});
  always
    @(posedge clk) begin
      reg220 <= ($unsigned($signed(reg119[(2'h3):(1'h0)])) && ((($signed(reg119) ?
          $unsigned(reg125) : $signed(wire219)) ^~ wire219[(4'h8):(3'h6)]) == reg122[(2'h2):(1'h1)]));
    end
  always
    @(posedge clk) begin
      if ({($signed(wire131) > (+$signed((reg122 ? reg122 : reg118)))),
          (|$unsigned((~|{reg119})))})
        begin
          reg221 <= $unsigned($signed(reg123[(3'h7):(1'h0)]));
          if ((8'hb7))
            begin
              reg222 <= (~(reg122[(3'h5):(2'h3)] <= {{$signed(reg125),
                      (+reg118)}}));
              reg223 <= ((&(&$unsigned(reg117[(3'h6):(3'h4)]))) >> {reg222});
            end
          else
            begin
              reg222 <= (~wire109[(4'ha):(3'h5)]);
              reg223 <= (|($unsigned({wire113[(1'h0):(1'h0)], wire112}) ?
                  $unsigned($unsigned(reg128[(2'h2):(1'h0)])) : $unsigned($signed((wire219 + wire108)))));
              reg224 <= $unsigned($unsigned(reg221[(1'h1):(1'h1)]));
              reg225 <= reg124[(2'h2):(1'h0)];
              reg226 <= ({(8'hab),
                  {(&$unsigned((8'ha8)))}} != wire108[(3'h5):(3'h5)]);
            end
        end
      else
        begin
          reg221 <= $signed((!$signed({(reg116 ? reg129 : (8'hba))})));
          reg222 <= (-(wire111[(2'h2):(2'h2)] - $signed(reg119)));
          reg223 <= {$unsigned((((-wire108) ?
                      $signed(reg117) : (reg127 <<< reg117)) ?
                  {$signed(reg226)} : reg115))};
          reg224 <= wire108;
          reg225 <= {reg117[(5'h12):(4'he)], reg122[(3'h5):(2'h3)]};
        end
      reg227 <= (+(~^({(^~wire112),
          (reg126 < reg115)} != ({reg118} << wire109[(4'h9):(3'h5)]))));
      reg228 <= {$unsigned((~^wire219[(2'h2):(1'h1)]))};
    end
  assign wire229 = reg123;
  always
    @(posedge clk) begin
      reg230 <= ((($unsigned($signed(reg124)) == wire108[(2'h2):(1'h0)]) <<< {(~|{wire114}),
          ((-wire132) >>> $signed(reg125))}) && $signed(reg121));
      if ((+($unsigned($unsigned(wire114)) ?
          ({(reg120 >= reg127)} <<< wire229[(4'he):(3'h5)]) : $signed($unsigned((reg119 ^ wire108))))))
        begin
          reg231 <= ($signed((~|wire219)) < (reg127 ?
              ((+{reg117, reg225}) ?
                  {wire229[(3'h7):(3'h4)]} : (8'hae)) : ((7'h40) ?
                  reg122 : $signed((reg126 ? reg119 : wire108)))));
          reg232 <= (|reg127);
          reg233 <= (reg126[(3'h6):(2'h2)] == reg117);
        end
      else
        begin
          reg231 <= reg122;
          reg232 <= $signed($unsigned({(~|(reg128 ? reg226 : wire111))}));
          reg233 <= $unsigned((~|((8'ha2) ?
              {(reg220 ? reg127 : reg225), $unsigned(reg129)} : ((wire112 ?
                      (7'h40) : reg115) ?
                  (reg127 ? (8'ha7) : reg123) : (-(8'hac))))));
          reg234 <= reg126[(4'hf):(3'h7)];
          reg235 <= wire108[(1'h0):(1'h0)];
        end
      reg236 <= wire131[(4'hc):(3'h4)];
    end
  assign wire237 = (reg233 ?
                       {wire131[(4'hd):(3'h5)],
                           $unsigned((^~(~&reg123)))} : (((|{reg236, (8'ha8)}) ?
                               (~reg119[(4'h9):(4'h9)]) : {$unsigned(reg129),
                                   (8'hb9)}) ?
                           $signed(reg228[(5'h10):(2'h2)]) : $unsigned((-$signed((8'hbc))))));
  assign wire238 = $unsigned(reg118[(2'h3):(2'h2)]);
  assign wire239 = {$unsigned((($signed(reg129) ?
                           (reg129 ? (8'haa) : reg225) : (reg226 ?
                               reg226 : reg235)) << $signed((reg225 ?
                           reg126 : reg120)))),
                       {reg224, $signed(($signed(wire112) ? reg118 : reg125))}};
  assign wire240 = $signed($signed(reg235));
endmodule

module module4_1
#( parameter param86 = ((({((7'h41) <= (8'ha6))} ? (|{(8'hbd), (8'hbd)}) : (8'hb3)) ? ((-((8'h9c) ? (7'h43) : (8'h9c))) && (-((8'h9e) ? (8'ha8) : (8'h9d)))) : (({(8'h9d)} >= ((8'haf) <= (8'haf))) ^~ ((8'ha9) | (~^(8'hb9))))) ? (~&((((8'hbe) ~^ (8'h9e)) ? (~(8'ha2)) : ((8'ha1) ? (8'hb7) : (8'ha6))) ? (((8'hb4) >>> (8'hbb)) <= (8'hb6)) : (((8'ha0) ? (8'h9c) : (7'h42)) ? {(8'ha7), (8'h9e)} : (&(8'haf))))) : ((^~(((8'ha4) + (8'hac)) ? ((8'haf) > (8'ha8)) : ((8'ha9) && (8'hbd)))) > ((~&(^~(8'hbf))) || (!{(7'h40), (8'ha9)}))))
, parameter param87 = (param86 ? ((8'ha2) ? {((!param86) > (param86 ? param86 : param86)), param86} : ((~(param86 + param86)) > ((param86 ? param86 : (8'h9c)) ? param86 : {(8'h9d), param86}))) : (((7'h41) || (param86 ? (+param86) : (param86 ^~ param86))) >= (((param86 > param86) + (param86 ? param86 : param86)) ? ((8'ha2) <<< (~&param86)) : ((~&param86) && {param86})))) )
(y, clk, wire8, wire7, wire6, wire5);
  output wire [(32'h135):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire8;
  input wire signed [(5'h14):(1'h0)] wire7;
  input wire signed [(3'h6):(1'h0)] wire6;
  input wire signed [(5'h14):(1'h0)] wire5;
  wire signed [(3'h5):(1'h0)] wire85;
  wire signed [(4'hf):(1'h0)] wire38;
  wire [(4'ha):(1'h0)] wire10;
  wire signed [(5'h12):(1'h0)] wire9;
  wire [(4'hd):(1'h0)] wire40;
  reg signed [(5'h15):(1'h0)] reg41 = (1'h0);
  reg [(2'h2):(1'h0)] reg42 = (1'h0);
  reg [(4'ha):(1'h0)] reg43 = (1'h0);
  reg [(4'hf):(1'h0)] reg44 = (1'h0);
  reg [(2'h2):(1'h0)] reg45 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg46 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg47 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg48 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg49 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg50 = (1'h0);
  reg [(5'h15):(1'h0)] reg51 = (1'h0);
  wire [(4'hc):(1'h0)] wire52;
  wire signed [(4'hc):(1'h0)] wire53;
  wire [(4'h8):(1'h0)] wire54;
  wire signed [(4'hd):(1'h0)] wire55;
  wire signed [(4'h9):(1'h0)] wire56;
  wire [(4'hd):(1'h0)] wire57;
  wire [(2'h2):(1'h0)] wire58;
  wire signed [(3'h6):(1'h0)] wire59;
  wire signed [(3'h7):(1'h0)] wire60;
  wire signed [(3'h6):(1'h0)] wire61;
  wire signed [(4'ha):(1'h0)] wire62;
  wire [(5'h10):(1'h0)] wire83;
  assign y = {wire85,
                 wire38,
                 wire10,
                 wire9,
                 wire40,
                 reg41,
                 reg42,
                 reg43,
                 reg44,
                 reg45,
                 reg46,
                 reg47,
                 reg48,
                 reg49,
                 reg50,
                 reg51,
                 wire52,
                 wire53,
                 wire54,
                 wire55,
                 wire56,
                 wire57,
                 wire58,
                 wire59,
                 wire60,
                 wire61,
                 wire62,
                 wire83,
                 (1'h0)};
  assign wire9 = wire8[(2'h2):(1'h1)];
  assign wire10 = $unsigned(wire5[(1'h0):(1'h0)]);
  module11_1 modinst39 (wire38, clk, wire6, wire7, wire9, wire8, wire5);
  assign wire40 = $unsigned({{{$unsigned((8'hb2)), (wire10 >= wire7)}},
                      ($signed((+wire8)) << {wire5, (wire8 == wire10)})});
  always
    @(posedge clk) begin
      reg41 <= ({$unsigned($unsigned((wire8 ? (8'ha6) : wire8))),
              (|$signed(wire7[(3'h6):(2'h2)]))} ?
          (wire40[(2'h3):(1'h0)] ?
              (~|$signed((wire10 ?
                  wire38 : (8'hba)))) : $signed(wire5)) : $unsigned(wire5));
      reg42 <= (8'ha9);
      reg43 <= ((reg42 ^~ $unsigned((~(7'h40)))) ?
          (wire7 ? wire7 : wire38) : $signed(reg41));
      if ({{wire10[(2'h3):(1'h1)]}})
        begin
          reg44 <= (($signed(((7'h42) ?
                  $unsigned(reg42) : (wire5 ^~ wire10))) >= wire6) ?
              $signed((+$unsigned((|wire40)))) : wire6[(2'h3):(2'h3)]);
          reg45 <= $unsigned(reg42[(2'h2):(1'h0)]);
          reg46 <= $unsigned((^~wire6[(3'h6):(1'h0)]));
          reg47 <= (&$signed($unsigned(wire40)));
        end
      else
        begin
          reg44 <= wire6[(3'h6):(3'h5)];
          if ($unsigned((!$unsigned((wire40[(2'h3):(1'h0)] ^~ {reg42})))))
            begin
              reg45 <= wire10[(4'h9):(3'h5)];
              reg46 <= (reg47[(3'h6):(3'h6)] == (-($unsigned((reg43 ?
                  reg42 : wire40)) || wire6[(3'h6):(3'h5)])));
              reg47 <= reg41[(2'h3):(1'h1)];
              reg48 <= ((^~$unsigned({reg42,
                  ((8'ha3) - wire9)})) - ($signed(reg46[(4'ha):(4'h9)]) < ((~wire6[(3'h4):(3'h4)]) * $signed((7'h44)))));
            end
          else
            begin
              reg45 <= ((~(((reg41 ?
                  wire9 : wire7) ^~ wire9) ^ wire10[(3'h4):(1'h1)])) == (&(({wire5} >>> $signed(wire8)) ?
                  ((~wire10) >= (reg42 & (8'ha5))) : $unsigned((reg45 ?
                      wire10 : reg48)))));
              reg46 <= (reg43 < (~&{wire6[(3'h4):(1'h0)],
                  wire5[(1'h1):(1'h1)]}));
              reg47 <= ({(((&reg47) - $signed((8'haa))) + wire7)} ?
                  (reg47[(2'h3):(2'h2)] ?
                      (wire38[(4'hd):(1'h0)] ^~ $signed((reg48 ~^ reg45))) : reg43[(1'h1):(1'h1)]) : reg45);
            end
          reg49 <= wire40;
          reg50 <= (+$signed(reg42[(1'h1):(1'h0)]));
        end
      reg51 <= $signed($signed(wire8));
    end
  assign wire52 = (!reg47[(2'h2):(1'h1)]);
  assign wire53 = {wire40[(2'h2):(1'h1)], wire10[(4'h8):(3'h4)]};
  assign wire54 = ($unsigned($unsigned(wire10[(2'h2):(1'h0)])) ?
                      (reg43 ?
                          (&wire52[(1'h1):(1'h0)]) : (reg43[(1'h1):(1'h0)] <= wire10)) : ($signed(reg51[(4'h9):(1'h1)]) ^~ ($unsigned(reg45[(2'h2):(2'h2)]) != ($signed(wire5) ?
                          $unsigned(wire10) : wire10[(3'h6):(1'h0)]))));
  assign wire55 = $unsigned(wire52[(4'h9):(3'h6)]);
  assign wire56 = {(wire7 ?
                          wire40[(2'h3):(1'h1)] : (((wire52 ?
                                  wire38 : (8'hbf)) <= wire38) ?
                              $signed(wire54[(2'h3):(1'h0)]) : $signed(((8'hb0) ?
                                  wire10 : wire9)))),
                      $signed(wire10)};
  assign wire57 = $unsigned((-(reg50 ?
                      reg43[(2'h2):(2'h2)] : $unsigned($signed(wire54)))));
  assign wire58 = $unsigned(reg48);
  assign wire59 = {({((|reg46) ? $unsigned(reg51) : reg49)} ?
                          ({(wire9 ? (8'haf) : reg45)} != ($unsigned(reg41) ?
                              {reg51} : (wire57 <<< (8'ha9)))) : $unsigned((^~reg47[(2'h2):(1'h0)]))),
                      (-reg45[(1'h0):(1'h0)])};
  assign wire60 = $signed((((((8'hb8) ? (8'ha7) : wire58) ?
                          ((8'had) <<< reg42) : $signed((8'ha8))) * (-wire54[(3'h4):(2'h3)])) ?
                      (~^reg49[(4'h8):(4'h8)]) : wire56[(4'h8):(3'h4)]));
  assign wire61 = $unsigned($signed(wire54));
  assign wire62 = $signed((!$signed((~^wire6[(1'h0):(1'h0)]))));
  module63_1 modinst84 (.wire68(wire6), .wire64(wire55), .wire67(reg49), .clk(clk), .y(wire83), .wire66(reg43), .wire65(wire40));
  assign wire85 = wire54[(4'h8):(3'h7)];
endmodule

module module63_1
#( parameter param81 = (({(~(|(8'hac))), (~|((8'hb1) ? (7'h41) : (8'ha5)))} != ((((8'hab) < (7'h44)) ? (+(8'h9d)) : ((8'hae) << (8'ha3))) ? (&((8'ha2) >= (7'h41))) : (|(~^(8'hb7))))) <<< (({((8'hba) ? (8'h9d) : (8'hb4))} ? (((8'hb9) + (8'ha4)) & (~(8'ha6))) : {(^(7'h41))}) == {(8'hbc), ((~&(8'ha4)) ? ((8'hac) ~^ (8'ha8)) : ((8'hb6) ? (8'hb4) : (8'h9c)))}))
, parameter param82 = {param81, ((param81 >> ((param81 ? param81 : (7'h40)) ? (param81 & param81) : (^~param81))) ? (~&((param81 >> param81) < {(8'hbe), param81})) : param81)} )
(y, clk, wire68, wire67, wire66, wire65, wire64);
  output wire [(32'h77):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h4):(1'h0)] wire68;
  input wire signed [(2'h2):(1'h0)] wire67;
  input wire [(4'ha):(1'h0)] wire66;
  input wire [(4'hd):(1'h0)] wire65;
  input wire signed [(4'hb):(1'h0)] wire64;
  wire signed [(5'h10):(1'h0)] wire80;
  wire [(4'hf):(1'h0)] wire79;
  wire signed [(4'h9):(1'h0)] wire78;
  reg [(3'h4):(1'h0)] reg77 = (1'h0);
  reg [(4'h9):(1'h0)] reg76 = (1'h0);
  reg [(3'h5):(1'h0)] reg75 = (1'h0);
  reg [(5'h15):(1'h0)] reg74 = (1'h0);
  reg signed [(4'he):(1'h0)] reg73 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire72;
  wire [(3'h5):(1'h0)] wire71;
  wire [(4'h8):(1'h0)] wire70;
  wire [(3'h7):(1'h0)] wire69;
  assign y = {wire80,
                 wire79,
                 wire78,
                 reg77,
                 reg76,
                 reg75,
                 reg74,
                 reg73,
                 wire72,
                 wire71,
                 wire70,
                 wire69,
                 (1'h0)};
  assign wire69 = wire65;
  assign wire70 = ((^~$signed((wire69 ? $signed(wire64) : wire64))) + wire68);
  assign wire71 = wire65;
  assign wire72 = (8'hbc);
  always
    @(posedge clk) begin
      if (wire68)
        begin
          if ((wire72[(1'h1):(1'h0)] ?
              (wire68 ?
                  {($unsigned(wire68) >= (wire70 ? wire68 : (8'h9c))),
                      {$unsigned((8'ha2))}} : {(-$signed(wire65))}) : $signed($signed(wire72))))
            begin
              reg73 <= wire67;
              reg74 <= $unsigned(($unsigned(wire72) ?
                  wire70[(3'h7):(1'h0)] : $unsigned($unsigned($signed((7'h44))))));
              reg75 <= $signed($unsigned((~({(7'h44), wire64} != (wire67 ?
                  wire64 : wire66)))));
              reg76 <= (|(8'had));
            end
          else
            begin
              reg73 <= ({$signed((^(+reg73))),
                      ((reg75 ?
                          (wire70 ^ wire70) : (wire72 ?
                              wire72 : reg73)) <= {(~reg75)})} ?
                  {$unsigned($unsigned(reg75)),
                      {((8'ha6) || (reg75 ?
                              wire72 : wire64))}} : ((8'hb4) && reg73[(1'h1):(1'h1)]));
              reg74 <= $signed(reg74[(5'h15):(3'h5)]);
            end
        end
      else
        begin
          if ($signed($unsigned(wire69[(3'h6):(3'h5)])))
            begin
              reg73 <= (+wire67);
              reg74 <= $signed(reg75[(2'h3):(1'h1)]);
              reg75 <= {((wire64[(1'h1):(1'h0)] ^ (8'h9d)) <<< wire72),
                  {(^~({wire72} ~^ reg73[(4'hc):(3'h5)])),
                      {reg73[(4'hd):(3'h4)], (+reg75)}}};
              reg76 <= wire66[(1'h0):(1'h0)];
            end
          else
            begin
              reg73 <= (~|wire65[(3'h6):(1'h1)]);
              reg74 <= wire64;
              reg75 <= $unsigned(((~&reg73) >= $signed(wire64)));
            end
          reg77 <= (wire64[(4'h9):(3'h6)] ^ reg76);
        end
    end
  assign wire78 = ($signed($signed(reg74[(1'h0):(1'h0)])) << $signed(reg75[(1'h1):(1'h1)]));
  assign wire79 = (-(^~(reg74 <<< wire66)));
  assign wire80 = {reg75, {wire64}};
endmodule

module module11_1  (y, clk, wire16, wire15, wire14, wire13, wire12);
  output wire [(32'h11f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire16;
  input wire [(2'h2):(1'h0)] wire15;
  input wire [(4'h9):(1'h0)] wire14;
  input wire [(5'h11):(1'h0)] wire13;
  input wire [(4'h9):(1'h0)] wire12;
  reg [(5'h10):(1'h0)] reg37 = (1'h0);
  reg [(4'he):(1'h0)] reg36 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire35;
  wire [(5'h11):(1'h0)] wire34;
  reg [(5'h12):(1'h0)] reg33 = (1'h0);
  reg [(4'h9):(1'h0)] reg32 = (1'h0);
  reg [(5'h15):(1'h0)] reg31 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg30 = (1'h0);
  reg [(5'h10):(1'h0)] reg29 = (1'h0);
  reg [(4'ha):(1'h0)] reg28 = (1'h0);
  reg [(5'h10):(1'h0)] reg27 = (1'h0);
  reg [(2'h3):(1'h0)] reg26 = (1'h0);
  reg [(4'h9):(1'h0)] reg25 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg24 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg23 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire22;
  wire [(5'h12):(1'h0)] wire21;
  reg signed [(2'h2):(1'h0)] reg20 = (1'h0);
  reg [(3'h7):(1'h0)] reg19 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg18 = (1'h0);
  wire [(4'h8):(1'h0)] wire17;
  assign y = {reg37,
                 reg36,
                 wire35,
                 wire34,
                 reg33,
                 reg32,
                 reg31,
                 reg30,
                 reg29,
                 reg28,
                 reg27,
                 reg26,
                 reg25,
                 reg24,
                 reg23,
                 wire22,
                 wire21,
                 reg20,
                 reg19,
                 reg18,
                 wire17,
                 (1'h0)};
  assign wire17 = ({wire13, {(|$unsigned(wire16))}} ~^ (wire12 ^~ (8'ha1)));
  always
    @(posedge clk) begin
      reg18 <= wire16;
      reg19 <= ((reg18 ? reg18 : wire17) ?
          $signed($unsigned($unsigned((wire13 ?
              wire13 : wire14)))) : $signed((-(^(~|wire14)))));
      reg20 <= wire13;
    end
  assign wire21 = ((wire16[(1'h0):(1'h0)] >>> ($signed((wire17 >>> reg19)) ^ (wire13 ?
                          {wire12} : $unsigned(wire16)))) ?
                      wire15[(1'h1):(1'h1)] : wire16[(3'h5):(3'h5)]);
  assign wire22 = wire15[(2'h2):(1'h0)];
  always
    @(posedge clk) begin
      reg23 <= ($signed($unsigned((|(reg20 & wire21)))) ?
          ((+$unsigned($signed(reg20))) ^ $unsigned({((8'haa) ^~ (7'h40)),
              (!reg19)})) : $unsigned($unsigned(((reg19 ?
              wire16 : wire15) < {wire13}))));
      reg24 <= (wire22 ?
          $signed(wire15[(1'h0):(1'h0)]) : wire17[(2'h3):(1'h0)]);
      if ({wire13[(4'he):(1'h1)], (wire16 && (8'hb1))})
        begin
          reg25 <= (((wire14 ?
                      ((8'ha7) < (|reg20)) : ($unsigned(wire15) ?
                          (reg19 ? wire15 : reg19) : wire22[(1'h1):(1'h0)])) ?
                  (wire14[(4'h9):(3'h4)] && {wire17}) : {$unsigned((wire17 ?
                          wire12 : wire15))}) ?
              ((wire22[(4'h9):(3'h7)] | $unsigned({reg19})) ?
                  $signed(((wire17 ?
                      wire22 : wire12) && (reg23 * wire22))) : {$signed($signed(wire21))}) : {(({wire12} - wire15[(2'h2):(1'h1)]) ^~ $signed((-reg20))),
                  reg18});
          reg26 <= wire15[(1'h1):(1'h0)];
          reg27 <= (reg25 - (|$signed($unsigned((wire22 >>> reg18)))));
          if ({($signed({{wire12, reg26},
                  wire12[(2'h3):(2'h3)]}) < wire22[(5'h11):(3'h6)])})
            begin
              reg28 <= wire13;
              reg29 <= ((wire21[(2'h3):(1'h0)] ?
                      wire22[(2'h3):(2'h3)] : reg28) ?
                  ($unsigned({$signed(reg26)}) <<< ($signed((wire17 ?
                          reg23 : wire14)) ?
                      ({reg18, wire15} ?
                          (wire15 ?
                              reg24 : reg18) : $signed((8'h9c))) : $signed($signed(reg18)))) : $signed(reg27[(4'ha):(1'h0)]));
              reg30 <= reg29[(1'h1):(1'h1)];
              reg31 <= $unsigned((reg19 ?
                  {$signed((+reg25)),
                      $unsigned((wire13 ?
                          wire17 : reg27))} : $signed((reg23[(4'h8):(1'h1)] <<< wire12))));
            end
          else
            begin
              reg28 <= $unsigned(($unsigned($unsigned($signed(reg25))) ?
                  $unsigned(((reg19 <<< (8'h9f)) ^ (-(7'h42)))) : reg26));
              reg29 <= $signed(((^((reg25 ^ reg26) ?
                  reg31[(3'h4):(1'h1)] : reg18)) ^~ ((-$signed(reg25)) ?
                  {$unsigned(wire21)} : wire17[(3'h7):(3'h6)])));
            end
        end
      else
        begin
          reg25 <= $unsigned($signed((reg19 ?
              {$unsigned((8'hb2))} : $unsigned($signed(wire14)))));
          reg26 <= (~^((wire21 ?
                  $unsigned({(8'h9d), wire22}) : $signed($unsigned(reg26))) ?
              wire12[(3'h5):(1'h1)] : ($unsigned((|wire16)) ?
                  $signed($signed((8'hbf))) : reg31[(2'h2):(1'h1)])));
        end
      reg32 <= $signed(($unsigned((~|wire22[(2'h2):(2'h2)])) & (^~$unsigned((wire17 ?
          (8'hb0) : reg26)))));
    end
  always
    @(posedge clk) begin
      reg33 <= ((~|$signed($signed($signed(wire12)))) ?
          (reg19[(2'h3):(2'h2)] ^~ (reg23[(1'h0):(1'h0)] ?
              reg20 : reg30)) : (wire22 ?
              $signed(((!reg28) ?
                  (reg18 || reg18) : (wire13 >> wire13))) : wire21[(5'h12):(3'h4)]));
    end
  assign wire34 = wire13;
  assign wire35 = $signed(reg27[(2'h2):(2'h2)]);
  always
    @(posedge clk) begin
      reg36 <= wire14;
      reg37 <= wire35[(5'h11):(3'h7)];
    end
endmodule

module module133_1  (y, clk, wire137, wire136, wire135, wire134);
  output wire [(32'h355):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire137;
  input wire [(5'h14):(1'h0)] wire136;
  input wire signed [(4'hd):(1'h0)] wire135;
  input wire [(4'h9):(1'h0)] wire134;
  wire signed [(3'h7):(1'h0)] wire216;
  wire signed [(4'ha):(1'h0)] wire215;
  reg signed [(4'h9):(1'h0)] reg214 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg213 = (1'h0);
  reg [(4'ha):(1'h0)] reg212 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg211 = (1'h0);
  reg [(5'h13):(1'h0)] reg210 = (1'h0);
  reg [(4'hd):(1'h0)] reg209 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg208 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg207 = (1'h0);
  reg [(5'h13):(1'h0)] reg206 = (1'h0);
  reg signed [(4'he):(1'h0)] reg205 = (1'h0);
  reg [(3'h5):(1'h0)] reg204 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg203 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg202 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg201 = (1'h0);
  reg [(5'h15):(1'h0)] reg200 = (1'h0);
  reg [(3'h6):(1'h0)] reg199 = (1'h0);
  reg [(2'h2):(1'h0)] reg198 = (1'h0);
  reg signed [(4'he):(1'h0)] reg197 = (1'h0);
  reg [(4'ha):(1'h0)] reg196 = (1'h0);
  reg [(4'hc):(1'h0)] reg195 = (1'h0);
  wire [(4'ha):(1'h0)] wire194;
  reg signed [(4'hb):(1'h0)] reg193 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg192 = (1'h0);
  reg [(4'h8):(1'h0)] reg191 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg190 = (1'h0);
  reg [(4'hb):(1'h0)] reg189 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg188 = (1'h0);
  reg [(3'h6):(1'h0)] reg187 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg186 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg185 = (1'h0);
  reg [(5'h11):(1'h0)] reg184 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg183 = (1'h0);
  reg [(3'h6):(1'h0)] reg182 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg181 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg180 = (1'h0);
  reg [(3'h4):(1'h0)] reg179 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire178;
  wire [(4'hd):(1'h0)] wire177;
  wire signed [(4'he):(1'h0)] wire176;
  wire signed [(4'hc):(1'h0)] wire175;
  wire [(4'ha):(1'h0)] wire174;
  reg signed [(3'h4):(1'h0)] reg173 = (1'h0);
  reg [(3'h6):(1'h0)] reg172 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg171 = (1'h0);
  reg [(2'h3):(1'h0)] reg170 = (1'h0);
  reg [(5'h10):(1'h0)] reg169 = (1'h0);
  reg [(5'h10):(1'h0)] reg168 = (1'h0);
  reg [(2'h3):(1'h0)] reg167 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg166 = (1'h0);
  reg [(5'h15):(1'h0)] reg165 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg164 = (1'h0);
  reg [(5'h15):(1'h0)] reg163 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg162 = (1'h0);
  reg [(5'h12):(1'h0)] reg161 = (1'h0);
  reg [(4'hc):(1'h0)] reg160 = (1'h0);
  reg [(2'h3):(1'h0)] reg159 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg158 = (1'h0);
  reg [(5'h12):(1'h0)] reg157 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg156 = (1'h0);
  reg [(5'h14):(1'h0)] reg155 = (1'h0);
  reg [(2'h3):(1'h0)] reg154 = (1'h0);
  reg [(4'hf):(1'h0)] reg153 = (1'h0);
  reg [(4'hf):(1'h0)] reg152 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg151 = (1'h0);
  reg [(4'hc):(1'h0)] reg150 = (1'h0);
  wire [(5'h10):(1'h0)] wire149;
  reg [(4'hf):(1'h0)] reg148 = (1'h0);
  reg [(5'h15):(1'h0)] reg147 = (1'h0);
  reg [(2'h3):(1'h0)] reg146 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg145 = (1'h0);
  wire [(3'h4):(1'h0)] wire144;
  wire [(2'h3):(1'h0)] wire143;
  wire [(3'h5):(1'h0)] wire142;
  wire [(5'h11):(1'h0)] wire141;
  wire [(2'h3):(1'h0)] wire140;
  wire [(5'h12):(1'h0)] wire139;
  wire [(2'h3):(1'h0)] wire138;
  assign y = {wire216,
                 wire215,
                 reg214,
                 reg213,
                 reg212,
                 reg211,
                 reg210,
                 reg209,
                 reg208,
                 reg207,
                 reg206,
                 reg205,
                 reg204,
                 reg203,
                 reg202,
                 reg201,
                 reg200,
                 reg199,
                 reg198,
                 reg197,
                 reg196,
                 reg195,
                 wire194,
                 reg193,
                 reg192,
                 reg191,
                 reg190,
                 reg189,
                 reg188,
                 reg187,
                 reg186,
                 reg185,
                 reg184,
                 reg183,
                 reg182,
                 reg181,
                 reg180,
                 reg179,
                 wire178,
                 wire177,
                 wire176,
                 wire175,
                 wire174,
                 reg173,
                 reg172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 wire149,
                 reg148,
                 reg147,
                 reg146,
                 reg145,
                 wire144,
                 wire143,
                 wire142,
                 wire141,
                 wire140,
                 wire139,
                 wire138,
                 (1'h0)};
  assign wire138 = wire136;
  assign wire139 = $signed(((((wire134 ? wire138 : wire135) != wire135) ?
                       $signed((~^wire138)) : $unsigned({wire134})) < (&(+$signed(wire134)))));
  assign wire140 = (wire137[(3'h5):(1'h0)] ?
                       wire136[(4'hb):(3'h7)] : (~&$signed(wire136[(4'he):(2'h2)])));
  assign wire141 = {wire140[(1'h1):(1'h1)]};
  assign wire142 = (~($unsigned((!$signed(wire138))) * wire137[(3'h5):(3'h4)]));
  assign wire143 = ((+((wire136[(5'h12):(4'h9)] ^~ wire139) ?
                           $signed(wire142[(2'h3):(2'h2)]) : (~^wire140[(2'h3):(1'h0)]))) ?
                       ((^wire140[(2'h3):(1'h0)]) ?
                           $unsigned(({wire134} - wire137[(1'h1):(1'h0)])) : wire137[(4'h9):(3'h4)]) : ($unsigned((-wire138)) < ((wire142 ?
                           wire138[(1'h0):(1'h0)] : $unsigned(wire137)) * ((~^(8'hb9)) ?
                           (wire139 == wire138) : $unsigned(wire135)))));
  assign wire144 = (&{$unsigned({{wire135, wire141}, (~&wire139)}), wire139});
  always
    @(posedge clk) begin
      reg145 <= $signed((7'h43));
      reg146 <= {$signed((-($signed(wire139) - wire139[(4'hb):(4'h8)]))),
          reg145[(2'h3):(2'h3)]};
      reg147 <= wire142[(2'h2):(2'h2)];
      reg148 <= ($unsigned((^~((wire134 ?
              wire140 : reg147) != $signed(wire140)))) ?
          ((((!wire138) ~^ (wire142 ? wire140 : (8'h9c))) ?
                  reg147 : $signed($unsigned(wire139))) ?
              (({wire134, wire143} * (wire134 < wire142)) ?
                  $unsigned($signed(reg146)) : $signed($signed(wire136))) : (($signed(wire134) < (wire138 ?
                      wire138 : wire136)) ?
                  $signed(wire134[(3'h4):(2'h2)]) : $unsigned((reg146 ?
                      wire141 : wire143)))) : wire135);
    end
  assign wire149 = wire138[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      reg150 <= (((8'hb8) && (8'h9c)) > ($signed(((wire137 || (8'hba)) >> (+(8'hb7)))) ?
          $signed(wire138) : $unsigned($signed($signed(reg147)))));
      if ((^~($unsigned(wire135) < ((+(|wire143)) && ($unsigned(reg146) >= {reg147,
          reg145})))))
        begin
          reg151 <= wire137[(4'h9):(2'h3)];
          if ({wire138[(1'h0):(1'h0)]})
            begin
              reg152 <= (|reg150);
              reg153 <= ({$unsigned({reg146[(2'h3):(2'h2)], $unsigned(reg147)}),
                      (8'ha2)} ?
                  $unsigned((reg152[(1'h0):(1'h0)] ?
                      wire144 : $unsigned((-wire135)))) : $unsigned(wire149));
            end
          else
            begin
              reg152 <= $unsigned((^reg151[(2'h2):(1'h1)]));
              reg153 <= (wire140[(1'h1):(1'h1)] ?
                  {$unsigned({(wire138 ? wire140 : wire136),
                          $unsigned(wire144)})} : $signed((((reg153 >> (8'hb2)) ?
                          {reg152, reg152} : wire149) ?
                      (^~$unsigned(wire138)) : (^$signed(wire142)))));
              reg154 <= ($signed($signed(((^~wire149) ?
                      wire143 : (^wire141)))) ?
                  reg146 : $unsigned((wire135 ?
                      wire149[(4'ha):(2'h3)] : wire139[(5'h12):(3'h7)])));
            end
          reg155 <= (!wire135[(3'h6):(3'h4)]);
          reg156 <= (|(($signed(wire142[(2'h3):(1'h1)]) ?
              wire142 : {(reg150 ? reg148 : wire137)}) & wire137));
        end
      else
        begin
          reg151 <= ((^(^(-(wire144 > wire143)))) == (wire137 ?
              wire141 : reg151));
          reg152 <= reg153;
          reg153 <= ((({$unsigned(wire140),
                  $signed((8'hab))} ^ $signed(wire138)) ^ (~{$unsigned(wire136)})) ?
              (7'h41) : (reg156[(1'h0):(1'h0)] ?
                  (-{wire140}) : $signed($signed((^reg153)))));
        end
      if (wire135)
        begin
          reg157 <= $unsigned($unsigned($unsigned($signed((~&reg147)))));
          if (((($unsigned((~|wire138)) ^ ($unsigned(reg157) >>> (reg155 ?
                  wire143 : reg155))) <= ((~(wire139 ?
                  wire135 : wire139)) >>> (wire144[(1'h1):(1'h1)] ?
                  (|(8'hac)) : wire142[(2'h2):(1'h1)]))) ?
              wire138 : $unsigned((((reg157 ? reg146 : wire138) + (~^wire141)) ?
                  ((8'hb1) ^ (reg157 || wire142)) : {wire135, reg148}))))
            begin
              reg158 <= $unsigned(reg151[(2'h3):(2'h3)]);
              reg159 <= ($unsigned({wire134[(3'h5):(2'h3)],
                      (~&wire139[(1'h1):(1'h1)])}) ?
                  $signed(reg156) : (wire142[(1'h1):(1'h1)] ?
                      $signed(wire141) : (~|($unsigned(wire134) ?
                          (^wire142) : ((8'h9f) ? wire136 : reg155)))));
              reg160 <= reg145[(3'h4):(2'h3)];
              reg161 <= (((wire144 ?
                      (~^(^~wire134)) : $signed((~wire134))) + (^~$signed(reg159))) ?
                  ($signed((~^reg154)) ?
                      $signed(reg154[(2'h3):(1'h0)]) : reg156) : ($unsigned(wire144) > wire143));
              reg162 <= reg147;
            end
          else
            begin
              reg158 <= $unsigned((~reg158));
            end
          reg163 <= wire143[(2'h3):(2'h2)];
          if (reg146)
            begin
              reg164 <= ($signed(($unsigned((wire144 ?
                      wire136 : (8'hae))) * $unsigned((reg145 ?
                      reg159 : (8'hba))))) ?
                  ((8'hb4) ?
                      wire135[(4'h8):(3'h6)] : ($signed((^reg160)) ?
                          (8'hbf) : $unsigned(wire143[(2'h3):(2'h2)]))) : ({$unsigned(reg155),
                      $signed($signed(reg151))} <<< wire139[(4'h9):(2'h2)]));
              reg165 <= (+$unsigned(reg151[(1'h0):(1'h0)]));
              reg166 <= $signed($signed(((+wire149) ?
                  wire144[(1'h1):(1'h1)] : $signed((~&wire137)))));
              reg167 <= (~($unsigned((8'hab)) >> (+reg148)));
              reg168 <= $signed($signed(((8'hb4) ?
                  ((wire142 ? wire137 : reg158) * $signed(reg153)) : (8'hb4))));
            end
          else
            begin
              reg164 <= ((8'hb5) ?
                  $signed({reg154[(2'h2):(2'h2)],
                      (wire142[(3'h5):(1'h0)] <<< (wire144 < reg164))}) : reg159);
              reg165 <= {((8'ha6) ? $unsigned($signed(reg152)) : (8'ha1))};
            end
          if (($unsigned((reg163 ?
              (wire135[(2'h3):(1'h0)] == reg165[(2'h2):(2'h2)]) : (~|{reg159,
                  (8'hb4)}))) == ($unsigned(wire142) == wire140)))
            begin
              reg169 <= (~&reg165);
              reg170 <= reg157;
            end
          else
            begin
              reg169 <= (+wire135);
              reg170 <= wire144;
              reg171 <= $signed({($signed($signed((7'h40))) ?
                      ((~|(8'ha7)) ?
                          (^reg162) : $unsigned(reg152)) : (8'ha0))});
              reg172 <= (+($unsigned((reg159[(2'h3):(2'h2)] ?
                  {reg152} : (~wire141))) > (($signed(reg166) ?
                  (~&wire144) : $signed(reg168)) & reg160)));
              reg173 <= wire134[(1'h0):(1'h0)];
            end
        end
      else
        begin
          reg157 <= reg152;
          reg158 <= {$unsigned($unsigned(reg168[(2'h3):(1'h0)])),
              (reg146 > $signed(((reg169 ?
                  wire141 : reg155) * (reg158 < (8'hbc)))))};
          if (wire136[(5'h14):(5'h13)])
            begin
              reg159 <= reg160[(3'h4):(2'h2)];
              reg160 <= (wire134[(1'h0):(1'h0)] ^ $signed($unsigned($unsigned((~^wire142)))));
            end
          else
            begin
              reg159 <= $signed($signed($signed((+reg166))));
              reg160 <= reg147;
              reg161 <= (((|$unsigned({(8'haa)})) ?
                      reg172[(1'h1):(1'h1)] : {(^reg170), reg164}) ?
                  ({{reg166[(4'hb):(3'h6)], reg145[(2'h2):(1'h0)]},
                      (-{reg162})} >>> reg156) : ((~$unsigned($unsigned(reg170))) ~^ $signed((~|$signed(reg162)))));
              reg162 <= $unsigned(reg172);
            end
          reg163 <= {{reg159, ((^~((8'hb9) ? reg166 : reg153)) ^ wire141)}};
          if ($unsigned(((reg148[(4'hc):(3'h5)] ?
              (reg167 > reg165[(4'ha):(3'h7)]) : wire142[(1'h1):(1'h0)]) * $signed($unsigned((reg170 ?
              reg158 : (8'ha8)))))))
            begin
              reg164 <= $signed((reg173 ?
                  (((reg145 ^ wire149) ?
                      (reg170 <= wire140) : (wire140 || (8'hbf))) * ((~wire136) | (8'hba))) : $unsigned(({reg166,
                          reg169} ?
                      $unsigned(wire134) : {reg162, reg162}))));
              reg165 <= (-((reg151 ?
                  reg156[(1'h1):(1'h1)] : $unsigned($signed(reg146))) & wire139));
              reg166 <= (8'ha1);
              reg167 <= ($signed(reg158[(1'h1):(1'h1)]) ?
                  wire135[(2'h2):(2'h2)] : $unsigned((&(^~((7'h44) >= (8'ha4))))));
            end
          else
            begin
              reg164 <= (($signed((&$signed((8'ha4)))) <= wire149[(1'h0):(1'h0)]) ?
                  $unsigned($unsigned(reg159)) : ($unsigned(wire144[(1'h0):(1'h0)]) && reg166));
              reg165 <= (&$unsigned(reg171));
              reg166 <= $signed($unsigned(({{wire140}} ? {wire141} : reg163)));
            end
        end
    end
  assign wire174 = reg167[(1'h1):(1'h0)];
  assign wire175 = wire139[(4'hd):(1'h1)];
  assign wire176 = (~^(((reg146[(1'h1):(1'h0)] ?
                           (!reg167) : ((8'haf) ? wire174 : reg146)) ?
                       wire138[(1'h0):(1'h0)] : $unsigned(reg153[(2'h2):(1'h0)])) ~^ reg166));
  assign wire177 = (8'hba);
  assign wire178 = wire142[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      if (($unsigned((^((^~reg167) <= reg162[(4'hd):(2'h2)]))) > {(wire176[(4'hb):(4'ha)] ?
              ($unsigned(reg150) <<< (reg171 ?
                  wire139 : (8'hae))) : (&$unsigned(wire175))),
          (wire149 ? (8'haf) : $unsigned(reg167[(2'h2):(1'h1)]))}))
        begin
          reg179 <= $signed($signed($unsigned($signed((reg169 ?
              reg168 : reg150)))));
          reg180 <= reg179[(1'h1):(1'h1)];
          if ($unsigned(((7'h40) << reg163[(5'h14):(4'h8)])))
            begin
              reg181 <= reg161;
            end
          else
            begin
              reg181 <= reg158[(5'h12):(5'h11)];
              reg182 <= reg171[(2'h2):(1'h0)];
              reg183 <= wire149;
              reg184 <= {(-(&(~&{wire175})))};
              reg185 <= {$unsigned((~$unsigned((wire141 - wire176)))),
                  $unsigned((reg165[(4'hc):(3'h4)] <= (!$signed(reg155))))};
            end
          reg186 <= $signed($unsigned(($signed(((8'hb8) || reg172)) + reg184)));
        end
      else
        begin
          if (((($signed((reg172 ? wire139 : reg162)) == {(reg185 ?
                          wire177 : (8'h9f))}) ?
                  $unsigned(((!reg152) ?
                      $signed(reg163) : $unsigned((8'hba)))) : reg148) ?
              ((8'ha5) & ({$signed(wire149),
                  $signed(reg160)} >= (((8'h9c) >>> reg170) ?
                  $signed(reg163) : ((8'haa) ?
                      reg170 : wire139)))) : $signed((((reg171 <= (8'ha4)) ?
                      $signed((8'ha4)) : (7'h43)) ?
                  {$unsigned((8'hb0)),
                      reg156} : ((reg157 != reg160) ~^ wire134[(3'h6):(1'h1)])))))
            begin
              reg179 <= $signed((wire139 ?
                  reg171 : {(reg180 ~^ $unsigned(reg153))}));
              reg180 <= $signed((&reg150));
              reg181 <= $unsigned(reg162);
            end
          else
            begin
              reg179 <= reg158;
              reg180 <= $signed($signed((~&((reg163 | (8'ha4)) ^~ $signed(reg161)))));
              reg181 <= (reg157 ? wire135 : $unsigned($signed(wire176)));
              reg182 <= (-(7'h40));
            end
          reg183 <= $unsigned($signed(reg173));
          reg184 <= (^{{(reg169 ? (reg155 >> reg179) : {reg145}),
                  (((8'h9f) ^~ reg148) ?
                      (reg156 ? reg186 : reg186) : (wire178 <<< reg165))},
              ($signed(reg146[(1'h0):(1'h0)]) ?
                  (~&(7'h41)) : $signed((reg150 <= reg154)))});
          reg185 <= reg182;
        end
      if (reg162)
        begin
          reg187 <= reg156[(1'h1):(1'h1)];
        end
      else
        begin
          reg187 <= (reg145 - (&wire175[(3'h7):(2'h2)]));
          reg188 <= (|$unsigned((reg145[(4'ha):(2'h3)] || (7'h42))));
          reg189 <= reg181;
          if ($unsigned(reg148[(4'ha):(4'h8)]))
            begin
              reg190 <= (&(({(reg157 ? reg188 : wire135)} ?
                  reg162[(1'h1):(1'h0)] : {(reg160 ?
                          wire174 : (8'ha4))}) ^~ reg180[(2'h2):(1'h1)]));
              reg191 <= ($unsigned(wire176) ?
                  $unsigned(reg183[(3'h4):(3'h4)]) : wire144);
            end
          else
            begin
              reg190 <= reg163;
            end
          reg192 <= wire137;
        end
    end
  always
    @(posedge clk) begin
      reg193 <= {((~^{wire134[(2'h3):(1'h0)], {reg167, wire138}}) ?
              $signed($signed($signed(reg169))) : (^$signed((wire137 << reg146)))),
          (^reg191[(3'h7):(1'h1)])};
    end
  assign wire194 = $unsigned($signed((-reg182)));
  always
    @(posedge clk) begin
      reg195 <= (~^reg152);
      if ({$unsigned(($signed((reg192 <= wire143)) >> ((wire174 ?
                  wire134 : (8'hbe)) ?
              (~^reg158) : $unsigned(reg158)))),
          reg165})
        begin
          reg196 <= (|(reg155 < reg185));
        end
      else
        begin
          reg196 <= (|($unsigned($unsigned(wire149)) ?
              ($unsigned(wire134) - (wire144 ?
                  $signed((8'hb6)) : (8'h9d))) : (7'h42)));
          reg197 <= {(&(~($unsigned((8'ha1)) ? $signed(wire137) : reg188)))};
        end
      reg198 <= $signed((!($signed($unsigned((7'h42))) ?
          (reg187[(1'h1):(1'h0)] * wire178) : wire194[(4'ha):(4'h8)])));
      reg199 <= {wire149};
      if (({$unsigned({(reg198 == reg166)})} ?
          (~^(((~|reg189) * $unsigned(wire177)) || ($unsigned(reg163) - (-reg184)))) : wire142))
        begin
          if ((-$signed($unsigned(((~&reg186) ? (reg173 + reg182) : reg150)))))
            begin
              reg200 <= reg162[(4'h8):(1'h0)];
              reg201 <= ($unsigned(reg168) == $signed(($signed((~&reg185)) == (reg163[(5'h13):(4'hf)] ?
                  $signed(reg159) : $unsigned(reg151)))));
              reg202 <= $signed((~reg183));
              reg203 <= (((wire142[(2'h3):(2'h2)] - wire140) ?
                  reg190[(1'h0):(1'h0)] : wire136) ^ reg201);
              reg204 <= (&{(&$unsigned((!reg198)))});
            end
          else
            begin
              reg200 <= (|{$signed((reg185 ?
                      $unsigned((8'hbb)) : $unsigned(reg189))),
                  ($unsigned($unsigned(reg185)) < $signed(wire177))});
            end
          if ((wire141 ~^ (^reg193)))
            begin
              reg205 <= $signed(wire177);
              reg206 <= $unsigned($signed(reg148[(3'h6):(3'h6)]));
              reg207 <= (~(reg181[(1'h0):(1'h0)] - $signed((+reg163[(4'hc):(3'h4)]))));
            end
          else
            begin
              reg205 <= reg206;
              reg206 <= wire136;
              reg207 <= (+reg157[(1'h0):(1'h0)]);
              reg208 <= (~&(!$signed(reg173[(3'h4):(1'h0)])));
            end
          if ($signed((~reg182[(3'h4):(1'h0)])))
            begin
              reg209 <= reg147;
              reg210 <= $signed(((8'ha5) || $signed((-$signed(reg205)))));
              reg211 <= ((((|$signed(wire137)) >= reg172[(3'h4):(2'h3)]) <<< $unsigned((&(reg173 ?
                  reg154 : reg156)))) <= reg199);
              reg212 <= (($unsigned($signed((reg158 == reg209))) ?
                  $signed((&(^reg204))) : (reg198[(1'h1):(1'h0)] ?
                      (reg201 ?
                          (reg171 == reg206) : (wire178 ?
                              (8'hbf) : (8'hac))) : (8'ha8))) - $unsigned($signed($signed($unsigned(reg184)))));
              reg213 <= $unsigned($unsigned(wire135));
            end
          else
            begin
              reg209 <= $unsigned(($unsigned(((reg209 & (8'ha6)) ?
                  $signed(reg161) : (~^reg213))) <<< (reg151 ?
                  reg168[(3'h5):(1'h1)] : $signed((reg211 ?
                      reg204 : reg197)))));
            end
          reg214 <= reg171[(2'h2):(1'h1)];
        end
      else
        begin
          reg200 <= $signed(($unsigned(wire135) ?
              ((!reg162) ?
                  $signed($unsigned((8'ha5))) : $unsigned((reg198 ?
                      reg179 : reg204))) : ($signed((wire175 >>> reg163)) ?
                  (reg153[(3'h4):(2'h3)] ? reg207 : (~^reg172)) : reg210)));
          if ($signed((wire194[(2'h3):(2'h3)] >= $signed(wire141))))
            begin
              reg201 <= {$unsigned(($unsigned((!reg171)) * {reg172}))};
              reg202 <= $signed(reg213);
              reg203 <= wire177;
              reg204 <= reg189[(4'h9):(1'h0)];
              reg205 <= {(+((wire174 ? $unsigned(wire139) : reg158) ?
                      $signed(wire149[(2'h2):(1'h0)]) : (-{reg170, reg170}))),
                  (((~|$signed(wire137)) < reg148[(3'h7):(1'h1)]) ?
                      $unsigned(((reg172 ^~ reg208) ?
                          reg189[(4'h9):(4'h9)] : $unsigned(reg168))) : $unsigned(((wire138 | wire149) ?
                          (&reg203) : $unsigned(reg206))))};
            end
          else
            begin
              reg201 <= {(8'hb7)};
            end
          reg206 <= $unsigned(((reg207[(2'h3):(2'h2)] >> ((reg210 ~^ reg160) ?
              $unsigned(reg173) : (reg164 ? reg192 : reg168))) ~^ {reg197,
              (wire140[(2'h2):(1'h1)] && (^reg205))}));
        end
    end
  assign wire215 = (reg173 <= (wire141[(4'hc):(1'h1)] ?
                       reg201 : ($signed($unsigned((8'h9d))) > reg151)));
  assign wire216 = (&{$signed($unsigned((reg200 ? reg164 : reg145)))});
endmodule