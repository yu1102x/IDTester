module top_1
#( parameter param270 = ({(8'h9c), ((((7'h40) ? (8'ha6) : (8'hb4)) >>> ((8'ha7) ? (8'hb0) : (8'ha0))) > {((8'ha0) ? (7'h42) : (8'ha4))})} ? (&({{(8'hae)}} + ((~|(8'ha0)) != ((8'ha4) >> (7'h40))))) : (((|((8'ha6) + (8'ha5))) <= (((8'hb0) ? (8'h9c) : (7'h44)) ? ((8'ha6) ? (8'hb0) : (8'hb4)) : (!(8'hb3)))) | ((~|((8'ha7) ? (8'hb0) : (8'h9d))) ? {((8'hbe) <<< (8'hbf)), ((8'ha8) ? (8'hb0) : (8'ha6))} : {(^(8'hb3)), (~&(8'ha6))}))) )
(y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'hc6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h13):(1'h0)] wire3;
  input wire [(5'h13):(1'h0)] wire2;
  input wire [(4'hc):(1'h0)] wire1;
  input wire [(4'ha):(1'h0)] wire0;
  wire [(4'ha):(1'h0)] wire269;
  wire signed [(5'h10):(1'h0)] wire268;
  wire signed [(4'hf):(1'h0)] wire112;
  wire [(5'h11):(1'h0)] wire4;
  wire [(4'h9):(1'h0)] wire251;
  wire signed [(4'hc):(1'h0)] wire253;
  wire signed [(5'h12):(1'h0)] wire254;
  wire signed [(3'h4):(1'h0)] wire255;
  wire [(3'h7):(1'h0)] wire256;
  wire signed [(4'h9):(1'h0)] wire258;
  wire signed [(2'h3):(1'h0)] wire259;
  wire [(3'h4):(1'h0)] wire260;
  wire signed [(5'h13):(1'h0)] wire261;
  wire [(5'h11):(1'h0)] wire262;
  wire [(4'ha):(1'h0)] wire263;
  wire [(4'h9):(1'h0)] wire264;
  wire [(5'h10):(1'h0)] wire265;
  wire [(2'h2):(1'h0)] wire266;
  assign y = {wire269,
                 wire268,
                 wire112,
                 wire4,
                 wire251,
                 wire253,
                 wire254,
                 wire255,
                 wire256,
                 wire258,
                 wire259,
                 wire260,
                 wire261,
                 wire262,
                 wire263,
                 wire264,
                 wire265,
                 wire266,
                 (1'h0)};
  assign wire4 = wire3[(1'h0):(1'h0)];
  module5_1 modinst113 (wire112, clk, wire0, wire3, wire4, wire2, wire1);
  module114_1 modinst252 (wire251, clk, wire1, wire2, wire4, wire112);
  assign wire253 = wire3;
  assign wire254 = wire251[(3'h7):(1'h0)];
  assign wire255 = ($unsigned(($signed((wire251 >>> wire253)) || $unsigned((~wire3)))) ?
                       ({wire0,
                           ($signed((8'ha7)) ^~ $unsigned(wire112))} & wire4) : $unsigned(($unsigned((wire112 != wire0)) - wire253[(4'hc):(1'h1)])));
  module37_1 modinst257 (.y(wire256), .wire41(wire253), .wire39(wire2), .wire40(wire4), .wire38(wire3), .clk(clk));
  assign wire258 = wire254[(1'h0):(1'h0)];
  assign wire259 = (&$signed($signed((!(wire253 ? (8'hb4) : wire2)))));
  assign wire260 = ($signed(wire258) >= $unsigned($unsigned((!wire253))));
  assign wire261 = $signed({(~&(8'hbf)), (~&wire259[(1'h0):(1'h0)])});
  assign wire262 = wire255;
  assign wire263 = wire258[(1'h1):(1'h0)];
  assign wire264 = wire4;
  assign wire265 = {(|wire2[(4'hd):(2'h3)])};
  module175_1 modinst267 (wire266, clk, wire0, wire2, wire265, wire251, wire254);
  assign wire268 = (($unsigned($signed({(8'ha8)})) << wire1) ?
                       wire112 : wire258);
  assign wire269 = (-((($unsigned((7'h41)) ?
                           $signed(wire4) : (wire258 < wire255)) > ((wire256 ?
                               wire254 : wire251) ?
                           $signed(wire253) : wire256)) ?
                       $signed($unsigned(wire258[(3'h7):(1'h1)])) : $unsigned((wire0 >>> (wire260 ?
                           (8'ha7) : (8'hb0))))));
endmodule

module module114_1  (y, clk, wire118, wire117, wire116, wire115);
  output wire [(32'h18d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire118;
  input wire [(3'h7):(1'h0)] wire117;
  input wire signed [(4'he):(1'h0)] wire116;
  input wire [(4'hf):(1'h0)] wire115;
  wire [(5'h12):(1'h0)] wire250;
  wire [(3'h4):(1'h0)] wire249;
  reg [(2'h3):(1'h0)] reg248 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg247 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg246 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg245 = (1'h0);
  reg [(4'hd):(1'h0)] reg244 = (1'h0);
  reg [(5'h12):(1'h0)] reg243 = (1'h0);
  wire [(4'h9):(1'h0)] wire242;
  wire signed [(3'h7):(1'h0)] wire241;
  reg signed [(4'h8):(1'h0)] reg240 = (1'h0);
  reg [(4'hd):(1'h0)] reg239 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg238 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg237 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire235;
  wire signed [(4'hd):(1'h0)] wire199;
  wire signed [(5'h14):(1'h0)] wire198;
  wire signed [(5'h10):(1'h0)] wire197;
  wire [(5'h11):(1'h0)] wire169;
  reg [(4'hd):(1'h0)] reg127 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg126 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg125 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg124 = (1'h0);
  reg [(5'h15):(1'h0)] reg123 = (1'h0);
  reg [(4'he):(1'h0)] reg122 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg121 = (1'h0);
  wire [(3'h4):(1'h0)] wire120;
  wire signed [(4'h9):(1'h0)] wire119;
  wire signed [(5'h15):(1'h0)] wire171;
  wire signed [(4'hf):(1'h0)] wire172;
  wire signed [(4'ha):(1'h0)] wire173;
  wire signed [(5'h12):(1'h0)] wire174;
  wire signed [(3'h4):(1'h0)] wire195;
  assign y = {wire250,
                 wire249,
                 reg248,
                 reg247,
                 reg246,
                 reg245,
                 reg244,
                 reg243,
                 wire242,
                 wire241,
                 reg240,
                 reg239,
                 reg238,
                 reg237,
                 wire235,
                 wire199,
                 wire198,
                 wire197,
                 wire169,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 reg121,
                 wire120,
                 wire119,
                 wire171,
                 wire172,
                 wire173,
                 wire174,
                 wire195,
                 (1'h0)};
  assign wire119 = ($signed($signed({((8'ha0) << wire116),
                       $unsigned((8'hba))})) | ((wire116 ?
                           wire117 : ($signed((8'haa)) <= (wire115 ?
                               wire116 : wire118))) ?
                       wire117[(2'h2):(1'h1)] : $unsigned(wire117)));
  assign wire120 = ({($signed((wire117 && wire118)) ?
                           (7'h42) : {$signed(wire115),
                               wire118})} ^~ $signed((($signed(wire117) ?
                           wire118[(1'h0):(1'h0)] : (wire119 & wire119)) ?
                       $signed(wire117) : wire119[(3'h7):(2'h3)])));
  always
    @(posedge clk) begin
      reg121 <= wire120[(1'h1):(1'h1)];
      reg122 <= wire117;
      if ($signed(wire115[(2'h2):(2'h2)]))
        begin
          if ({wire119,
              {{($signed(wire118) != (wire117 ? reg122 : wire119)),
                      ((wire117 ? wire118 : wire117) <= ((7'h41) * reg122))}}})
            begin
              reg123 <= {$unsigned({$unsigned(wire117[(2'h2):(1'h0)])})};
              reg124 <= $signed(reg121[(2'h3):(2'h2)]);
            end
          else
            begin
              reg123 <= reg124[(4'ha):(4'h9)];
            end
          reg125 <= wire116;
        end
      else
        begin
          if ((wire119[(1'h0):(1'h0)] ?
              $unsigned(wire118[(1'h1):(1'h0)]) : ((8'ha7) & $signed((+reg125[(3'h5):(1'h1)])))))
            begin
              reg123 <= wire117[(2'h2):(1'h1)];
              reg124 <= {(~$signed((&(wire120 > (8'hae))))),
                  (|((wire120 >> $unsigned((8'haf))) ?
                      {(8'h9d), {wire120}} : $signed((~^reg124))))};
              reg125 <= $signed($unsigned($unsigned((!$signed(wire116)))));
              reg126 <= (!(|$unsigned(reg122[(4'h9):(3'h4)])));
              reg127 <= wire117[(3'h4):(1'h0)];
            end
          else
            begin
              reg123 <= (|(-(($unsigned(wire119) ^~ $unsigned(reg126)) == reg126)));
              reg124 <= ((8'h9d) && (&(^~$unsigned((^wire116)))));
              reg125 <= reg125;
              reg126 <= reg121;
              reg127 <= (+reg124[(4'h8):(2'h3)]);
            end
        end
    end
  module128_1 modinst170 (.clk(clk), .y(wire169), .wire132(reg125), .wire131(reg123), .wire133(reg127), .wire130(wire115), .wire129(wire116));
  assign wire171 = wire120;
  assign wire172 = (reg126[(1'h1):(1'h1)] ?
                       $unsigned($unsigned(reg124[(4'hc):(4'ha)])) : $unsigned(({$signed(wire119)} ?
                           wire171[(5'h13):(1'h0)] : wire117[(2'h3):(1'h1)])));
  assign wire173 = $signed((-reg125));
  assign wire174 = $signed($signed($unsigned((wire169 > (8'haa)))));
  module175_1 modinst196 (wire195, clk, reg127, wire116, wire171, reg123, wire174);
  assign wire197 = reg125;
  assign wire198 = (8'ha4);
  assign wire199 = ($unsigned(reg124[(4'hb):(4'hb)]) - $signed({{(wire169 ?
                               (8'hb6) : wire171),
                           reg121},
                       ((|reg125) ?
                           (reg121 ? reg124 : wire115) : $unsigned(wire117))}));
  module200_1 modinst236 (.wire203(reg121), .y(wire235), .wire204(wire115), .wire201(wire118), .clk(clk), .wire202(wire116));
  always
    @(posedge clk) begin
      reg237 <= $unsigned(wire195[(1'h0):(1'h0)]);
      reg238 <= $unsigned(reg237[(2'h2):(1'h0)]);
      reg239 <= (reg237 ?
          ((|((wire117 ? reg121 : reg126) ?
              (~^wire198) : wire119)) & (reg124[(3'h7):(3'h7)] ~^ (8'ha7))) : reg123[(4'hf):(4'h9)]);
      reg240 <= reg237;
    end
  assign wire241 = (wire235[(1'h0):(1'h0)] ?
                       wire116[(4'he):(4'ha)] : reg126[(4'hc):(2'h3)]);
  assign wire242 = $signed((wire171 ?
                       (wire169[(4'ha):(4'h8)] ?
                           (^(wire120 * wire174)) : ({wire173} & (reg127 ~^ wire235))) : ((wire115 ?
                           (^~wire116) : reg122[(1'h0):(1'h0)]) + wire118[(3'h5):(2'h3)])));
  always
    @(posedge clk) begin
      reg243 <= wire174[(4'hc):(3'h6)];
      if (wire118)
        begin
          reg244 <= (((reg127 ?
                  wire119 : wire198) & $unsigned($unsigned(((8'hb3) ?
                  wire116 : reg240)))) ?
              reg239[(3'h4):(1'h1)] : ((^~wire118) ?
                  (|$unsigned((^reg121))) : $signed(wire197[(2'h2):(2'h2)])));
          reg245 <= (($signed(((~wire198) ?
              {(8'hbe)} : $unsigned(wire195))) ^ $signed(reg122[(3'h6):(3'h4)])) - {(&wire242[(3'h5):(1'h0)]),
              ($unsigned($unsigned(reg122)) >> (wire242[(3'h7):(1'h0)] << $unsigned(wire115)))});
          reg246 <= ((^{$unsigned(((8'hb2) ? wire120 : (8'h9d))),
                  (~|(+wire235))}) ?
              (|(({wire241, wire169} ?
                  (reg244 != reg122) : $signed(reg123)) != (!(8'had)))) : {wire195[(3'h4):(2'h2)],
                  $unsigned({(+wire117), (reg237 <= wire174)})});
          reg247 <= ({($unsigned(((8'ha8) <= reg246)) & (reg122[(4'he):(4'ha)] ?
                      (reg244 ^~ reg123) : {wire172})),
                  ((((8'ha0) > reg126) ~^ (wire173 ?
                      wire173 : wire198)) != $signed($unsigned(reg127)))} ?
              ($unsigned($unsigned({wire198,
                  reg124})) <<< (wire242[(4'h8):(2'h3)] << wire195)) : (+(+$signed((reg124 ~^ (8'ha8))))));
          reg248 <= (^{$signed($unsigned((reg123 | wire171)))});
        end
      else
        begin
          reg244 <= (8'hb5);
          reg245 <= (((~^$signed($signed(wire171))) ^ (~|((8'hb9) ~^ reg246))) ?
              $unsigned(reg123[(4'h8):(1'h0)]) : reg248[(1'h0):(1'h0)]);
        end
    end
  assign wire249 = reg243[(4'hb):(4'h8)];
  assign wire250 = $signed(reg248[(2'h3):(2'h3)]);
endmodule

module module5_1  (y, clk, wire10, wire9, wire8, wire7, wire6);
  output wire [(32'hfb):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire10;
  input wire [(5'h13):(1'h0)] wire9;
  input wire signed [(5'h11):(1'h0)] wire8;
  input wire [(4'hd):(1'h0)] wire7;
  input wire signed [(4'ha):(1'h0)] wire6;
  wire [(4'hc):(1'h0)] wire111;
  reg [(4'hf):(1'h0)] reg110 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg109 = (1'h0);
  reg [(3'h5):(1'h0)] reg108 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg107 = (1'h0);
  reg [(3'h4):(1'h0)] reg106 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg105 = (1'h0);
  wire [(4'h9):(1'h0)] wire104;
  wire [(4'h9):(1'h0)] wire103;
  wire [(5'h13):(1'h0)] wire102;
  reg signed [(4'he):(1'h0)] reg101 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg100 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire99;
  wire signed [(5'h11):(1'h0)] wire97;
  wire signed [(5'h11):(1'h0)] wire36;
  wire [(3'h5):(1'h0)] wire35;
  wire [(4'he):(1'h0)] wire34;
  wire [(5'h13):(1'h0)] wire32;
  wire signed [(5'h12):(1'h0)] wire12;
  wire [(5'h15):(1'h0)] wire11;
  assign y = {wire111,
                 reg110,
                 reg109,
                 reg108,
                 reg107,
                 reg106,
                 reg105,
                 wire104,
                 wire103,
                 wire102,
                 reg101,
                 reg100,
                 wire99,
                 wire97,
                 wire36,
                 wire35,
                 wire34,
                 wire32,
                 wire12,
                 wire11,
                 (1'h0)};
  assign wire11 = wire8;
  assign wire12 = $signed($unsigned($signed((~(wire11 ? (8'hbf) : wire11)))));
  module13_1 modinst33 (.clk(clk), .wire16(wire11), .wire17(wire10), .wire15(wire7), .wire14(wire12), .y(wire32));
  assign wire34 = $signed(wire10);
  assign wire35 = ($signed($signed((~wire9[(4'hc):(4'ha)]))) ?
                      (wire10[(3'h6):(1'h0)] & ($unsigned(((8'hac) ?
                              wire12 : wire32)) ?
                          ($unsigned(wire10) != wire34[(1'h0):(1'h0)]) : ((wire8 ?
                                  wire7 : wire6) ?
                              (wire32 ?
                                  (7'h44) : wire7) : $unsigned(wire34)))) : {wire12[(1'h0):(1'h0)],
                          wire10});
  assign wire36 = (({(wire10[(3'h5):(3'h5)] ?
                              (wire10 ? wire35 : wire10) : $signed(wire11)),
                          ((!wire12) > (|wire11))} ?
                      wire6 : $signed((8'ha6))) * (|$unsigned(((wire6 ?
                      wire9 : wire12) + (wire9 ^~ wire11)))));
  module37_1 modinst98 (wire97, clk, wire34, wire8, wire32, wire36);
  assign wire99 = (8'hac);
  always
    @(posedge clk) begin
      reg100 <= wire12;
      reg101 <= wire99;
    end
  assign wire102 = $unsigned(reg101[(4'hd):(4'h9)]);
  assign wire103 = wire8;
  assign wire104 = wire97;
  always
    @(posedge clk) begin
      reg105 <= $signed(wire8[(3'h6):(3'h4)]);
      if ((8'ha5))
        begin
          reg106 <= $signed((!(-(wire35 ? reg105 : (~^wire103)))));
          reg107 <= ((+$unsigned(wire34[(3'h4):(2'h3)])) & (8'h9f));
        end
      else
        begin
          reg106 <= ((-{(~^wire102[(4'h8):(4'h8)]),
              ((wire12 * wire99) ?
                  {wire8,
                      wire36} : reg101[(4'hc):(3'h6)])}) ~^ wire7[(4'h8):(1'h0)]);
          reg107 <= wire34;
        end
      reg108 <= $signed((8'hb4));
      reg109 <= (({$signed((+wire32))} + wire7[(3'h6):(2'h3)]) >= $signed($signed($signed((wire103 ?
          reg105 : wire12)))));
      reg110 <= reg101[(2'h3):(2'h3)];
    end
  assign wire111 = reg105;
endmodule

module module37_1  (y, clk, wire41, wire40, wire39, wire38);
  output wire [(32'h2ab):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire41;
  input wire [(5'h11):(1'h0)] wire40;
  input wire signed [(5'h13):(1'h0)] wire39;
  input wire signed [(5'h11):(1'h0)] wire38;
  wire signed [(3'h4):(1'h0)] wire96;
  wire [(4'hf):(1'h0)] wire95;
  wire signed [(5'h11):(1'h0)] wire94;
  wire signed [(5'h14):(1'h0)] wire93;
  wire [(5'h12):(1'h0)] wire92;
  reg [(5'h15):(1'h0)] reg91 = (1'h0);
  reg [(5'h11):(1'h0)] reg90 = (1'h0);
  reg [(5'h11):(1'h0)] reg89 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg88 = (1'h0);
  reg [(5'h15):(1'h0)] reg87 = (1'h0);
  reg [(5'h12):(1'h0)] reg86 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg85 = (1'h0);
  reg [(5'h11):(1'h0)] reg84 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg83 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg82 = (1'h0);
  reg [(4'ha):(1'h0)] reg81 = (1'h0);
  reg [(5'h11):(1'h0)] reg80 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg79 = (1'h0);
  reg [(4'ha):(1'h0)] reg78 = (1'h0);
  reg [(5'h13):(1'h0)] reg77 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg76 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg75 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg74 = (1'h0);
  reg [(4'hb):(1'h0)] reg73 = (1'h0);
  reg [(4'h8):(1'h0)] reg72 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg71 = (1'h0);
  reg [(3'h5):(1'h0)] reg70 = (1'h0);
  wire [(5'h13):(1'h0)] wire69;
  wire [(5'h15):(1'h0)] wire68;
  wire signed [(3'h7):(1'h0)] wire67;
  wire signed [(4'ha):(1'h0)] wire66;
  wire [(4'ha):(1'h0)] wire65;
  wire signed [(5'h12):(1'h0)] wire64;
  reg signed [(3'h6):(1'h0)] reg63 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg62 = (1'h0);
  reg [(5'h12):(1'h0)] reg61 = (1'h0);
  reg [(5'h10):(1'h0)] reg60 = (1'h0);
  reg [(4'h9):(1'h0)] reg59 = (1'h0);
  reg [(4'ha):(1'h0)] reg58 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg57 = (1'h0);
  reg [(5'h13):(1'h0)] reg56 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg55 = (1'h0);
  reg [(3'h6):(1'h0)] reg54 = (1'h0);
  reg [(5'h11):(1'h0)] reg53 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg52 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg51 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg50 = (1'h0);
  reg [(4'he):(1'h0)] reg49 = (1'h0);
  wire [(3'h7):(1'h0)] wire48;
  wire [(4'ha):(1'h0)] wire47;
  wire [(2'h2):(1'h0)] wire46;
  wire signed [(4'hc):(1'h0)] wire45;
  wire [(5'h10):(1'h0)] wire44;
  wire signed [(3'h7):(1'h0)] wire43;
  wire signed [(5'h14):(1'h0)] wire42;
  assign y = {wire96,
                 wire95,
                 wire94,
                 wire93,
                 wire92,
                 reg91,
                 reg90,
                 reg89,
                 reg88,
                 reg87,
                 reg86,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 reg80,
                 reg79,
                 reg78,
                 reg77,
                 reg76,
                 reg75,
                 reg74,
                 reg73,
                 reg72,
                 reg71,
                 reg70,
                 wire69,
                 wire68,
                 wire67,
                 wire66,
                 wire65,
                 wire64,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 reg55,
                 reg54,
                 reg53,
                 reg52,
                 reg51,
                 reg50,
                 reg49,
                 wire48,
                 wire47,
                 wire46,
                 wire45,
                 wire44,
                 wire43,
                 wire42,
                 (1'h0)};
  assign wire42 = $unsigned(($signed($signed($unsigned(wire39))) & ($signed($signed(wire41)) != ((^~wire41) <<< wire39))));
  assign wire43 = wire40[(4'hf):(3'h6)];
  assign wire44 = $signed((($unsigned((!wire38)) >= ((!wire39) ^~ (wire43 ^ (8'ha0)))) ?
                      $unsigned((wire41[(2'h3):(1'h0)] != {wire40})) : (($unsigned(wire40) ?
                              (wire41 ? wire43 : wire43) : $unsigned(wire39)) ?
                          ((+wire41) ?
                              wire38[(4'hd):(3'h5)] : $signed((8'h9e))) : ($unsigned(wire42) || $signed(wire40)))));
  assign wire45 = $unsigned(wire39[(3'h4):(3'h4)]);
  assign wire46 = $signed({($signed({wire40}) <= (~^$unsigned(wire44)))});
  assign wire47 = wire45[(4'hb):(4'ha)];
  assign wire48 = $signed({(!((wire39 ? wire39 : wire46) ^~ $signed(wire38))),
                      ($unsigned({wire47}) | wire47[(3'h4):(1'h1)])});
  always
    @(posedge clk) begin
      if (wire46)
        begin
          reg49 <= (wire42 ?
              wire38 : ((8'had) ?
                  {(wire45[(4'hb):(3'h5)] ?
                          (wire39 ? wire41 : (8'haf)) : $unsigned(wire44)),
                      {{wire46, wire48},
                          wire41[(3'h5):(2'h2)]}} : (^wire48[(1'h0):(1'h0)])));
          reg50 <= wire38;
          reg51 <= (8'ha3);
          if (({reg51[(4'hf):(4'hd)], wire47} ?
              $unsigned((-{$signed(wire40), wire48[(2'h2):(1'h0)]})) : wire46))
            begin
              reg52 <= (wire44 ^~ $unsigned(wire44[(4'hd):(3'h7)]));
              reg53 <= wire48[(1'h1):(1'h1)];
              reg54 <= (~(({(-wire38)} & $unsigned($signed(wire48))) | (~wire40)));
            end
          else
            begin
              reg52 <= (~&(wire47[(4'h9):(1'h0)] ?
                  $signed(((wire44 ? reg51 : reg49) ?
                      (wire43 ?
                          (8'hb0) : wire39) : (wire45 | wire39))) : ((~(wire42 * wire41)) ?
                      (~&(reg52 ? reg49 : reg52)) : wire44[(1'h1):(1'h1)])));
              reg53 <= wire38[(4'hc):(4'h9)];
              reg54 <= (-$unsigned((~$signed($signed(reg52)))));
            end
          reg55 <= {($unsigned(wire47) ?
                  ($signed($signed(reg53)) ?
                      wire38 : reg50[(1'h0):(1'h0)]) : ((+{wire47}) + $signed(((8'h9f) ?
                      wire41 : wire44)))),
              (($unsigned((~|reg54)) <= (wire38 ?
                      $signed(reg52) : (reg50 ? reg52 : reg51))) ?
                  {((~&(7'h42)) ? {wire39} : {reg52})} : (&(-reg51)))};
        end
      else
        begin
          reg49 <= ((wire44 ?
                  (({reg51} & $signed(wire47)) <<< wire44[(4'hd):(4'ha)]) : wire47) ?
              $signed(reg51) : $signed(($unsigned({reg54}) >> {$unsigned((8'hba))})));
        end
      reg56 <= $signed($unsigned(((wire40 ^~ (8'hab)) ?
          reg50[(1'h1):(1'h1)] : wire46[(1'h0):(1'h0)])));
      if ($signed((-$unsigned({$signed(reg50), (8'hb7)}))))
        begin
          reg57 <= wire42;
        end
      else
        begin
          reg57 <= $signed((~{($unsigned(reg54) <<< $unsigned(wire41))}));
          if ((&((reg49[(4'hb):(4'hb)] ? (-(~^wire46)) : reg54) ?
              ({(~^wire40), wire45[(4'h8):(1'h1)]} ?
                  $signed((wire47 >> (8'hae))) : (!$signed((8'ha3)))) : (8'h9e))))
            begin
              reg58 <= ($unsigned({(7'h43)}) ?
                  (^{(8'hb3), (~^$signed(reg53))}) : wire44);
              reg59 <= (+(!reg49[(2'h3):(2'h2)]));
              reg60 <= $unsigned((reg51 ^ (($signed(wire38) >>> $signed(wire44)) + (~|{reg58}))));
              reg61 <= $unsigned(((^$signed((reg54 ? wire39 : reg52))) ?
                  reg57[(1'h0):(1'h0)] : (&wire44[(1'h0):(1'h0)])));
              reg62 <= {reg50, wire43[(3'h7):(1'h0)]};
            end
          else
            begin
              reg58 <= reg52;
              reg59 <= reg59;
              reg60 <= (reg50[(2'h3):(2'h3)] ? wire48 : reg61[(3'h5):(1'h1)]);
              reg61 <= ({wire47, $signed($unsigned(wire47))} ?
                  ((reg49[(3'h6):(1'h0)] - (reg59 ?
                      wire39 : $unsigned(reg49))) <= ($signed(wire45) ?
                      $signed(((8'hb2) | reg57)) : $unsigned(reg53[(4'hf):(3'h4)]))) : {(8'ha3)});
              reg62 <= ({(&reg54)} ?
                  $unsigned($signed(((reg49 ? reg60 : wire47) ?
                      ((8'h9e) ~^ reg57) : (reg62 ?
                          wire42 : reg51)))) : $signed(wire45));
            end
        end
      reg63 <= wire39[(5'h12):(3'h4)];
    end
  assign wire64 = (~wire41[(2'h3):(1'h1)]);
  assign wire65 = (wire44[(4'hc):(4'h9)] <<< $signed(wire46));
  assign wire66 = wire38[(4'h9):(3'h7)];
  assign wire67 = $signed((^(reg49 ?
                      $unsigned(wire44[(1'h1):(1'h1)]) : reg55[(2'h2):(1'h1)])));
  assign wire68 = (8'hbf);
  assign wire69 = ({reg53[(5'h10):(3'h6)],
                          (reg62 >>> $unsigned((wire41 ? wire47 : reg59)))} ?
                      ($signed($signed(reg50)) ?
                          ((!wire38) ^ ($unsigned(reg59) ^ $unsigned(reg59))) : reg50) : reg60);
  always
    @(posedge clk) begin
      reg70 <= ($unsigned({{(reg52 - reg51)},
          ((reg57 != wire41) ?
              reg56 : $unsigned((8'h9f)))}) >>> (wire69[(3'h4):(3'h4)] > ((+$unsigned(wire64)) | ((wire45 ^ wire43) ?
          $unsigned(reg63) : {wire66}))));
      reg71 <= ($signed((-$signed(reg49[(4'hb):(2'h3)]))) && (^~reg52));
      reg72 <= $unsigned({$signed((((8'had) ? (8'ha8) : wire47) ?
              wire46[(2'h2):(1'h1)] : {wire42, reg62}))});
      reg73 <= reg70[(1'h1):(1'h1)];
      reg74 <= {reg71, reg50};
    end
  always
    @(posedge clk) begin
      reg75 <= {{(~|{(|reg61)})}};
      reg76 <= ($unsigned($signed(wire69[(5'h10):(1'h0)])) ?
          (({$unsigned((8'ha8))} ?
              reg75[(2'h2):(1'h0)] : $signed(wire40[(4'hf):(3'h6)])) != (-$signed(wire45[(1'h1):(1'h0)]))) : reg63[(2'h3):(2'h2)]);
      if ((wire66[(3'h7):(3'h6)] ?
          (wire42[(2'h2):(2'h2)] * {((reg50 ?
                  reg63 : reg75) || $unsigned(wire67)),
              reg59}) : reg56))
        begin
          if ({{(~^(8'hb5))}, ((reg70 | $signed(reg61)) ^~ reg53)})
            begin
              reg77 <= $signed((8'hbd));
              reg78 <= wire48[(2'h2):(1'h0)];
              reg79 <= reg55;
            end
          else
            begin
              reg77 <= (-$unsigned($signed($unsigned(reg50))));
              reg78 <= reg77;
            end
        end
      else
        begin
          reg77 <= $signed(((reg79 ? reg54[(2'h2):(1'h1)] : {$signed(wire39)}) ?
              reg62[(1'h0):(1'h0)] : $signed($unsigned($unsigned((7'h44))))));
          reg78 <= reg56;
          reg79 <= (|($unsigned($signed((wire69 ?
              wire68 : reg61))) & reg58[(1'h1):(1'h1)]));
          reg80 <= (($unsigned($unsigned((&reg61))) ^~ ($signed(wire43[(2'h2):(1'h0)]) ~^ $signed((reg59 - reg77)))) + reg50);
          if ((!((((wire40 ?
                  reg78 : wire43) ~^ (reg49 - wire43)) < reg74[(2'h3):(1'h1)]) ?
              (wire48 ^ reg71[(2'h3):(1'h0)]) : (reg52[(3'h4):(3'h4)] && ($unsigned(reg55) ?
                  (reg71 < reg49) : $unsigned((8'hac)))))))
            begin
              reg81 <= reg58;
              reg82 <= ((wire45[(4'h8):(3'h5)] >= $unsigned((^~$unsigned((8'hb0))))) > $signed((reg73[(1'h0):(1'h0)] ?
                  $unsigned((&wire69)) : $unsigned(wire40[(4'h9):(2'h2)]))));
              reg83 <= {$unsigned($unsigned((~(wire45 ? reg81 : reg51))))};
              reg84 <= (($signed($signed((wire40 ? (8'h9e) : wire64))) ?
                      reg79 : {(7'h44), reg73[(4'hb):(2'h2)]}) ?
                  $unsigned(reg56[(5'h10):(4'he)]) : (!($unsigned(wire40) ?
                      {(~^reg72),
                          (reg73 ?
                              wire66 : reg70)} : (reg73 != (reg57 * wire67)))));
              reg85 <= (+reg72[(3'h6):(1'h1)]);
            end
          else
            begin
              reg81 <= ((|$unsigned((~^(reg78 + reg74)))) ?
                  wire44[(3'h7):(3'h5)] : reg60);
              reg82 <= {reg50};
            end
        end
      reg86 <= (|((^~($unsigned(reg76) ? (~^reg60) : (reg54 + reg78))) ?
          reg83[(2'h2):(1'h1)] : reg60[(4'hc):(1'h0)]));
      if ($unsigned((($signed(reg77[(1'h0):(1'h0)]) + reg63[(1'h0):(1'h0)]) ?
          (!$unsigned(wire46[(1'h0):(1'h0)])) : reg57[(1'h1):(1'h0)])))
        begin
          if (wire38)
            begin
              reg87 <= ((&reg49) ?
                  reg63 : ($signed($signed((!wire68))) ?
                      (-$unsigned($signed(reg49))) : $signed(((^reg81) ?
                          {reg49} : $signed((8'ha7))))));
            end
          else
            begin
              reg87 <= reg62[(2'h2):(1'h0)];
            end
          reg88 <= $unsigned($unsigned($unsigned((reg83[(2'h2):(1'h0)] + {wire44}))));
          reg89 <= $signed(($signed({(wire66 - (8'hb0)), $unsigned((8'hb3))}) ?
              $unsigned(((reg79 ?
                  wire45 : reg84) == $unsigned(reg63))) : $unsigned((reg61[(4'hd):(4'hc)] + $signed(wire47)))));
          reg90 <= (reg52 ? (8'ha8) : wire41[(2'h3):(2'h2)]);
          reg91 <= $unsigned((wire47[(1'h0):(1'h0)] ?
              $unsigned(((reg62 ~^ reg89) ?
                  (wire39 ?
                      reg60 : (8'ha6)) : reg80)) : $unsigned(wire66[(4'h9):(4'h9)])));
        end
      else
        begin
          if (({wire45,
              $signed({$signed(reg54),
                  (reg61 ?
                      reg91 : reg89)})} ^~ ((((wire41 * wire42) > wire68) << wire65) ?
              reg76 : wire67[(3'h7):(3'h4)])))
            begin
              reg87 <= ((~^$signed((wire65 - $signed(reg72)))) ?
                  (^~$unsigned($unsigned($unsigned((8'ha9))))) : (~&wire45));
              reg88 <= reg53[(4'hd):(2'h3)];
              reg89 <= (+((reg76 ?
                      $unsigned({reg84, (8'h9e)}) : (|{reg57, wire48})) ?
                  $signed($signed((+reg59))) : (reg61 ?
                      (^~$unsigned(reg85)) : $unsigned((!reg71)))));
              reg90 <= ((^$signed((reg74 || (reg78 * (8'hbb))))) ?
                  ((!$signed((reg78 + reg58))) ?
                      wire45 : $signed((8'ha7))) : reg53[(3'h6):(1'h0)]);
            end
          else
            begin
              reg87 <= wire40;
              reg88 <= wire48[(3'h4):(2'h3)];
              reg89 <= reg57[(1'h1):(1'h1)];
            end
        end
    end
  assign wire92 = (8'ha2);
  assign wire93 = {({$unsigned((wire92 > (8'ha0))),
                          $unsigned($signed((8'hae)))} && {$signed((reg71 != wire65))}),
                      $signed({$signed((reg52 ? wire39 : wire66))})};
  assign wire94 = (8'hb1);
  assign wire95 = reg76[(2'h3):(2'h2)];
  assign wire96 = reg73;
endmodule

module module13_1
#( parameter param30 = (({({(8'haf), (8'hb9)} < {(8'hb4), (8'ha8)})} ? ((~|(|(8'haf))) ? (((8'hba) ? (8'hb3) : (8'hb5)) ? ((8'h9d) * (8'haa)) : (^(8'hb7))) : ({(8'h9d)} ? ((8'hbf) ? (8'hb0) : (8'h9d)) : (+(8'hb7)))) : ((((8'hba) ? (8'ha9) : (8'ha9)) | (8'ha2)) != (((8'hbf) ? (8'hb8) : (8'hbf)) ^~ ((8'hab) ? (8'h9d) : (8'haf))))) ? {(((^~(7'h43)) ? (-(7'h43)) : ((8'ha7) >> (8'hbf))) ? {(~^(7'h43)), ((8'hb9) ? (8'haa) : (8'hac))} : (((8'hb7) == (8'hbe)) ? ((8'hbc) ? (7'h43) : (8'h9d)) : ((8'ha7) ? (8'hb0) : (8'h9f)))), (~^(&(~(8'h9e))))} : (!(&(-((8'hbb) ? (8'hbc) : (8'hb9))))))
, parameter param31 = ((param30 && (&(7'h42))) && (8'hbf)) )
(y, clk, wire17, wire16, wire15, wire14);
  output wire [(32'h7c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire17;
  input wire [(5'h15):(1'h0)] wire16;
  input wire signed [(4'hd):(1'h0)] wire15;
  input wire [(5'h12):(1'h0)] wire14;
  wire signed [(3'h7):(1'h0)] wire29;
  wire [(5'h11):(1'h0)] wire28;
  wire [(3'h4):(1'h0)] wire27;
  wire signed [(4'hd):(1'h0)] wire26;
  wire signed [(2'h3):(1'h0)] wire25;
  wire signed [(2'h3):(1'h0)] wire24;
  wire [(3'h5):(1'h0)] wire23;
  wire [(3'h7):(1'h0)] wire22;
  wire signed [(5'h11):(1'h0)] wire21;
  wire signed [(5'h11):(1'h0)] wire20;
  wire signed [(4'hf):(1'h0)] wire19;
  wire [(4'hf):(1'h0)] wire18;
  assign y = {wire29,
                 wire28,
                 wire27,
                 wire26,
                 wire25,
                 wire24,
                 wire23,
                 wire22,
                 wire21,
                 wire20,
                 wire19,
                 wire18,
                 (1'h0)};
  assign wire18 = (wire16 ?
                      ((^$unsigned(wire15[(3'h6):(3'h5)])) <<< (wire14[(4'he):(1'h0)] < $signed((wire16 ?
                          wire15 : wire14)))) : (~|($signed((wire17 ?
                          wire17 : wire16)) ~^ (~^(8'hb3)))));
  assign wire19 = $signed((wire14 ? wire15 : wire16[(3'h7):(2'h2)]));
  assign wire20 = (wire17[(4'h9):(2'h2)] ?
                      (wire18[(4'h9):(1'h0)] <<< {((wire15 == (8'ha0)) ?
                              $signed(wire19) : wire17)}) : ($signed(wire15[(4'h9):(4'h8)]) >= ($signed(((7'h44) ?
                          wire18 : wire16)) * ($signed((8'ha5)) ?
                          wire17 : wire15[(4'h8):(3'h4)]))));
  assign wire21 = wire18;
  assign wire22 = wire18[(4'hf):(2'h2)];
  assign wire23 = wire16[(3'h4):(1'h0)];
  assign wire24 = $signed($signed(wire23));
  assign wire25 = wire16[(5'h12):(1'h1)];
  assign wire26 = (!$signed($signed((8'had))));
  assign wire27 = (wire22[(2'h2):(1'h0)] <= $signed($unsigned($unsigned($signed(wire25)))));
  assign wire28 = (wire17 <<< $signed((~^wire15[(2'h3):(2'h3)])));
  assign wire29 = (-(+(($unsigned(wire25) >>> $unsigned(wire25)) ?
                      {wire18[(1'h0):(1'h0)]} : wire20[(3'h4):(1'h1)])));
endmodule

module module200_1
#( parameter param233 = (((-{(^~(7'h41))}) || (-(~^((7'h40) ^ (8'hb4))))) >> ((({(8'hb6)} ? {(8'hb5), (8'ha7)} : (^(7'h42))) & ({(8'had)} ~^ ((7'h44) ? (7'h44) : (8'hb3)))) ? (!(((8'ha7) * (8'ha0)) ? {(7'h44)} : (~(8'hab)))) : ((~(^(8'h9f))) ? {(&(8'h9e))} : {{(8'ha2), (8'ha6)}})))
, parameter param234 = (&param233) )
(y, clk, wire204, wire203, wire202, wire201);
  output wire [(32'hff):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire204;
  input wire signed [(2'h2):(1'h0)] wire203;
  input wire [(4'he):(1'h0)] wire202;
  input wire signed [(4'hc):(1'h0)] wire201;
  wire signed [(4'h9):(1'h0)] wire232;
  wire [(3'h6):(1'h0)] wire231;
  wire signed [(4'ha):(1'h0)] wire230;
  wire signed [(3'h7):(1'h0)] wire229;
  wire [(4'he):(1'h0)] wire228;
  wire signed [(4'h9):(1'h0)] wire227;
  wire signed [(4'ha):(1'h0)] wire226;
  wire signed [(3'h6):(1'h0)] wire225;
  wire signed [(4'h9):(1'h0)] wire224;
  wire [(4'h8):(1'h0)] wire223;
  reg signed [(3'h7):(1'h0)] reg222 = (1'h0);
  reg [(2'h2):(1'h0)] reg221 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg220 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg219 = (1'h0);
  reg [(4'hd):(1'h0)] reg218 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg217 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg216 = (1'h0);
  reg [(3'h6):(1'h0)] reg215 = (1'h0);
  reg signed [(4'he):(1'h0)] reg214 = (1'h0);
  reg [(3'h4):(1'h0)] reg213 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg212 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg211 = (1'h0);
  reg [(4'ha):(1'h0)] reg210 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg209 = (1'h0);
  reg [(3'h4):(1'h0)] reg208 = (1'h0);
  wire [(3'h5):(1'h0)] wire207;
  wire [(5'h11):(1'h0)] wire206;
  wire signed [(4'hf):(1'h0)] wire205;
  assign y = {wire232,
                 wire231,
                 wire230,
                 wire229,
                 wire228,
                 wire227,
                 wire226,
                 wire225,
                 wire224,
                 wire223,
                 reg222,
                 reg221,
                 reg220,
                 reg219,
                 reg218,
                 reg217,
                 reg216,
                 reg215,
                 reg214,
                 reg213,
                 reg212,
                 reg211,
                 reg210,
                 reg209,
                 reg208,
                 wire207,
                 wire206,
                 wire205,
                 (1'h0)};
  assign wire205 = $signed((wire204 ?
                       (^$unsigned((~|wire201))) : (~&$signed($unsigned(wire202)))));
  assign wire206 = ($signed(((~|(|(8'hb3))) && wire205)) && {(wire205[(2'h3):(2'h3)] ?
                           $unsigned($signed(wire205)) : $unsigned({(8'ha2),
                               wire204}))});
  assign wire207 = $unsigned((-((~|wire202) ^~ ($unsigned((8'haf)) ?
                       $signed(wire205) : ((8'ha8) ^~ (8'hb4))))));
  always
    @(posedge clk) begin
      if ((8'hb8))
        begin
          if ((8'hb8))
            begin
              reg208 <= $signed($unsigned($unsigned(wire203)));
              reg209 <= wire205;
              reg210 <= (|$signed({(8'hb9)}));
              reg211 <= $signed(((~|((wire201 ? wire202 : wire204) ?
                      wire203 : $signed(wire206))) ?
                  reg210 : reg209[(1'h0):(1'h0)]));
            end
          else
            begin
              reg208 <= (~&reg210);
              reg209 <= wire201[(1'h1):(1'h0)];
              reg210 <= (|((&reg208) > ($unsigned((^reg208)) & $unsigned($signed(reg208)))));
              reg211 <= ((~wire204[(1'h0):(1'h0)]) >>> ((~$unsigned(wire204)) << ((+(reg211 ?
                      wire205 : (8'h9e))) ?
                  $unsigned((wire206 * reg208)) : $unsigned((reg210 ?
                      reg209 : wire207)))));
            end
          reg212 <= ($signed(($unsigned(wire204[(2'h3):(2'h2)]) >>> wire206[(2'h3):(2'h2)])) >= $unsigned(wire204[(2'h3):(2'h2)]));
          reg213 <= reg210[(4'ha):(3'h4)];
          reg214 <= $unsigned($signed((~|wire201[(3'h5):(1'h0)])));
          if (wire202)
            begin
              reg215 <= (&wire205[(1'h1):(1'h0)]);
            end
          else
            begin
              reg215 <= $unsigned($unsigned(({$signed(wire202),
                  (wire201 ?
                      wire205 : wire202)} ^~ $unsigned(reg209[(3'h7):(3'h5)]))));
            end
        end
      else
        begin
          reg208 <= $signed({$signed(((^wire201) && {reg214}))});
          reg209 <= (wire201 && reg210[(3'h7):(2'h2)]);
          if (wire201)
            begin
              reg210 <= reg208;
              reg211 <= $signed(reg210[(2'h2):(1'h0)]);
              reg212 <= $unsigned((reg209[(1'h0):(1'h0)] ^~ $unsigned((reg214 ?
                  ((8'hb1) ? (7'h43) : wire207) : $signed(wire203)))));
              reg213 <= wire205[(4'hc):(1'h0)];
              reg214 <= {((wire201 <<< reg211) ?
                      reg212[(3'h5):(2'h2)] : $signed($signed(((8'ha2) ?
                          reg215 : reg214)))),
                  ((((wire202 == wire204) < (~reg211)) ?
                      $signed((reg213 ?
                          reg214 : reg213)) : $signed({wire206})) ~^ reg209[(4'h9):(3'h4)])};
            end
          else
            begin
              reg210 <= $unsigned(($unsigned($signed((reg209 | reg208))) ?
                  (reg213 ?
                      wire205[(3'h7):(3'h5)] : (~&$unsigned(reg211))) : (!(8'hb4))));
              reg211 <= wire205;
              reg212 <= $unsigned({(8'h9d)});
              reg213 <= $signed($signed((&{{(8'ha6), reg214}, (!wire206)})));
              reg214 <= ($signed((+wire206[(3'h7):(3'h5)])) ?
                  (wire202[(3'h4):(1'h0)] + $signed(((~^reg212) ?
                      $signed(reg213) : $signed((8'hb9))))) : $unsigned((~&((~^wire202) & (reg208 ?
                      wire206 : wire201)))));
            end
        end
      reg216 <= ($unsigned((($unsigned(wire207) ?
              $signed(reg212) : (&(8'hab))) ^~ ((wire205 ? reg215 : reg211) ?
              reg208 : $signed(reg213)))) ?
          (~|wire201) : (reg211[(3'h5):(2'h2)] ?
              reg214 : reg213[(2'h3):(2'h3)]));
      if ((|$unsigned(wire205[(4'h8):(3'h6)])))
        begin
          reg217 <= wire201;
          reg218 <= {wire205};
        end
      else
        begin
          reg217 <= ((8'ha9) ?
              (((~(reg218 ? reg211 : wire205)) ?
                      ({reg208} - {reg215}) : (7'h40)) ?
                  $unsigned($unsigned($unsigned(wire206))) : $signed((~^reg208))) : $unsigned((wire201[(1'h0):(1'h0)] * (~reg210))));
          reg218 <= {$unsigned((~^reg217))};
          reg219 <= wire202;
          reg220 <= wire207;
        end
      reg221 <= wire205;
      reg222 <= wire207;
    end
  assign wire223 = (reg218 << $signed(reg218[(2'h3):(1'h1)]));
  assign wire224 = reg212;
  assign wire225 = (&$unsigned($unsigned(((~&reg213) ?
                       reg208[(2'h3):(1'h1)] : (wire223 << reg214)))));
  assign wire226 = ((7'h40) && ((($unsigned(reg222) ?
                           reg218 : $unsigned(reg219)) >= $unsigned((7'h44))) ?
                       (wire206 >>> wire223) : (~^$signed((reg219 + reg209)))));
  assign wire227 = wire224;
  assign wire228 = {($unsigned($unsigned(reg222[(2'h2):(1'h1)])) == reg217[(5'h11):(2'h3)])};
  assign wire229 = (^~reg216);
  assign wire230 = reg209;
  assign wire231 = reg208[(2'h3):(2'h3)];
  assign wire232 = {wire228};
endmodule

module module175_1
#(parameter param194 = (-((|(&(|(8'haf)))) ^~ (^~(^{(8'hba)})))))
(y, clk, wire180, wire179, wire178, wire177, wire176);
  output wire [(32'hc2):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h3):(1'h0)] wire180;
  input wire signed [(2'h2):(1'h0)] wire179;
  input wire [(5'h10):(1'h0)] wire178;
  input wire [(3'h6):(1'h0)] wire177;
  input wire [(5'h12):(1'h0)] wire176;
  wire signed [(5'h11):(1'h0)] wire193;
  wire signed [(5'h15):(1'h0)] wire192;
  wire [(5'h12):(1'h0)] wire191;
  wire signed [(4'hf):(1'h0)] wire190;
  wire signed [(4'hd):(1'h0)] wire189;
  wire [(4'hf):(1'h0)] wire188;
  reg signed [(3'h5):(1'h0)] reg187 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg186 = (1'h0);
  reg [(4'he):(1'h0)] reg185 = (1'h0);
  reg [(5'h13):(1'h0)] reg184 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg183 = (1'h0);
  wire [(5'h11):(1'h0)] wire182;
  wire [(5'h15):(1'h0)] wire181;
  assign y = {wire193,
                 wire192,
                 wire191,
                 wire190,
                 wire189,
                 wire188,
                 reg187,
                 reg186,
                 reg185,
                 reg184,
                 reg183,
                 wire182,
                 wire181,
                 (1'h0)};
  assign wire181 = ({((-$unsigned(wire178)) ?
                           ({wire176} ?
                               (wire176 ?
                                   wire177 : (8'hb8)) : (wire178 != wire180)) : (wire178[(4'hc):(3'h4)] >>> (~wire179)))} | wire179[(1'h0):(1'h0)]);
  assign wire182 = wire181[(3'h6):(3'h4)];
  always
    @(posedge clk) begin
      reg183 <= $signed(((($unsigned(wire182) ?
              wire180[(1'h0):(1'h0)] : (&wire181)) ?
          wire180 : (wire176 ?
              wire176 : {wire176})) >= ($unsigned((wire178 || wire180)) ?
          (~|wire176) : {$signed(wire176), (-wire179)})));
      reg184 <= (-(&$unsigned(($signed(wire176) ?
          $signed(wire177) : (|wire178)))));
      reg185 <= ({{$signed(wire178), reg184[(4'hc):(2'h3)]},
              $unsigned($signed($unsigned((8'hb4))))} ?
          (8'hbb) : $unsigned($unsigned({(wire179 ? wire181 : reg184)})));
      reg186 <= (^~$signed(wire181[(4'hd):(4'ha)]));
      reg187 <= ((^~reg184[(4'ha):(3'h5)]) ?
          reg186[(1'h1):(1'h1)] : wire179[(2'h2):(1'h1)]);
    end
  assign wire188 = (($signed((|(wire178 ? reg184 : wire176))) ?
                           ((&wire182[(3'h6):(3'h4)]) ?
                               wire182[(3'h7):(2'h2)] : ({reg187} ?
                                   (reg187 ?
                                       reg184 : wire179) : (reg186 & wire176))) : {wire178[(3'h7):(2'h3)]}) ?
                       $unsigned($unsigned($unsigned(reg186))) : ($signed({$unsigned(wire177)}) ?
                           (&reg183[(1'h1):(1'h0)]) : $signed((reg187[(2'h3):(2'h2)] ?
                               ((8'hbb) ?
                                   (7'h40) : (8'ha9)) : (wire182 >>> (8'h9f))))));
  assign wire189 = ((^(&($unsigned(wire180) ?
                       wire177[(3'h4):(3'h4)] : {wire177}))) ~^ ((^{{(8'h9d)},
                       $signed(reg184)}) && (~|(wire188[(4'hf):(3'h6)] ?
                       (reg184 ^ reg187) : (wire188 ? wire177 : (8'ha7))))));
  assign wire190 = wire180[(1'h0):(1'h0)];
  assign wire191 = $unsigned(wire188);
  assign wire192 = reg187;
  assign wire193 = {$unsigned((($signed((8'ha9)) < $signed(wire179)) ?
                           $unsigned(reg183) : $signed((wire188 | wire176))))};
endmodule

module module128_1  (y, clk, wire133, wire132, wire131, wire130, wire129);
  output wire [(32'h1d5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire133;
  input wire signed [(3'h6):(1'h0)] wire132;
  input wire signed [(4'hc):(1'h0)] wire131;
  input wire signed [(4'hf):(1'h0)] wire130;
  input wire [(3'h6):(1'h0)] wire129;
  wire signed [(4'ha):(1'h0)] wire168;
  wire signed [(4'h9):(1'h0)] wire167;
  wire signed [(4'hf):(1'h0)] wire166;
  wire signed [(5'h12):(1'h0)] wire165;
  wire signed [(3'h6):(1'h0)] wire164;
  wire signed [(5'h13):(1'h0)] wire163;
  reg [(3'h5):(1'h0)] reg162 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg161 = (1'h0);
  reg [(5'h12):(1'h0)] reg160 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg159 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg158 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg157 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg156 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg155 = (1'h0);
  reg [(4'ha):(1'h0)] reg154 = (1'h0);
  reg [(3'h5):(1'h0)] reg153 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg152 = (1'h0);
  reg [(4'ha):(1'h0)] reg151 = (1'h0);
  reg [(4'h9):(1'h0)] reg150 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire149;
  wire signed [(4'ha):(1'h0)] wire148;
  reg signed [(4'he):(1'h0)] reg147 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg146 = (1'h0);
  reg [(5'h12):(1'h0)] reg145 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg144 = (1'h0);
  reg [(2'h3):(1'h0)] reg143 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg142 = (1'h0);
  reg [(2'h2):(1'h0)] reg141 = (1'h0);
  reg signed [(4'he):(1'h0)] reg140 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg139 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire138;
  reg [(5'h11):(1'h0)] reg137 = (1'h0);
  reg [(4'hd):(1'h0)] reg136 = (1'h0);
  wire [(2'h2):(1'h0)] wire135;
  wire [(5'h10):(1'h0)] wire134;
  assign y = {wire168,
                 wire167,
                 wire166,
                 wire165,
                 wire164,
                 wire163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 wire149,
                 wire148,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 reg143,
                 reg142,
                 reg141,
                 reg140,
                 reg139,
                 wire138,
                 reg137,
                 reg136,
                 wire135,
                 wire134,
                 (1'h0)};
  assign wire134 = $unsigned(wire130);
  assign wire135 = (((($unsigned(wire133) + wire131) == ($unsigned(wire133) ?
                               (+wire133) : (^(8'ha6)))) ?
                           (^(wire130[(1'h0):(1'h0)] ~^ wire133[(4'h8):(4'h8)])) : wire131[(4'ha):(1'h0)]) ?
                       (wire134 ?
                           wire129 : wire132[(3'h6):(1'h1)]) : $signed($unsigned(wire130[(2'h3):(2'h2)])));
  always
    @(posedge clk) begin
      reg136 <= wire130;
      reg137 <= wire133;
    end
  assign wire138 = wire135;
  always
    @(posedge clk) begin
      reg139 <= wire135[(1'h0):(1'h0)];
      if ((&wire129))
        begin
          reg140 <= $signed(wire134);
          reg141 <= (reg137[(5'h10):(3'h5)] ? wire132 : wire135);
          reg142 <= wire135;
          reg143 <= $signed(((+$signed((reg139 ? (8'hbf) : reg140))) ?
              (-$signed(wire133[(4'hd):(4'h9)])) : (reg139 ?
                  reg136[(3'h5):(1'h1)] : wire131)));
        end
      else
        begin
          if ({$signed($unsigned((-wire129[(2'h3):(2'h3)])))})
            begin
              reg140 <= (($signed({(reg139 - wire135),
                  $unsigned((8'ha3))}) != {(~wire132[(2'h2):(1'h1)])}) > (($signed($unsigned(reg140)) ?
                      (&(reg136 ^ wire132)) : ((reg143 ?
                          (7'h41) : reg139) ^~ wire138)) ?
                  $unsigned($unsigned($signed(wire130))) : (reg141[(1'h0):(1'h0)] ?
                      ($signed((8'h9e)) ?
                          reg140 : $signed((8'ha0))) : $unsigned((wire131 | wire130)))));
              reg141 <= (8'hb4);
              reg142 <= $signed(wire129);
              reg143 <= (|reg137[(4'ha):(3'h5)]);
              reg144 <= reg143;
            end
          else
            begin
              reg140 <= $signed((+$unsigned($signed($signed(wire135)))));
              reg141 <= (reg139 ? reg137 : (wire133[(1'h1):(1'h1)] * reg141));
              reg142 <= wire131;
            end
        end
      reg145 <= $unsigned((~^$signed(((!(8'ha1)) - (~&wire134)))));
      reg146 <= ((wire134[(3'h5):(3'h5)] >>> reg141[(1'h1):(1'h1)]) ~^ $unsigned($unsigned(reg145)));
      reg147 <= $signed($unsigned({wire133[(3'h4):(2'h2)],
          $unsigned({(7'h40), wire138})}));
    end
  assign wire148 = (|wire129);
  assign wire149 = wire131[(1'h1):(1'h1)];
  always
    @(posedge clk) begin
      reg150 <= ((~|{({reg137, (8'hb7)} ^~ (!wire131)),
              (reg139[(3'h4):(1'h0)] == (wire130 || (8'hbe)))}) ?
          wire132 : wire129);
      reg151 <= wire135;
      if ($unsigned((reg143[(2'h3):(1'h0)] ?
          (+$unsigned($unsigned(reg136))) : wire131)))
        begin
          if (({((^~{wire135, reg147}) ?
                      {$unsigned((8'ha7))} : (reg145 ?
                          reg151[(2'h3):(2'h3)] : {reg141, reg143}))} ?
              ((~&reg146[(3'h6):(3'h5)]) ?
                  $signed(wire129[(1'h0):(1'h0)]) : $signed($unsigned(wire130[(4'h9):(3'h5)]))) : (wire133[(4'hd):(4'h9)] ?
                  (^$unsigned(((8'h9e) * reg145))) : {$signed((reg144 || reg150)),
                      (+$signed(reg145))})))
            begin
              reg152 <= (wire132[(3'h6):(3'h6)] >>> ($unsigned($unsigned(wire134[(4'hc):(1'h0)])) && (((reg140 ?
                  reg143 : reg137) >>> reg143[(1'h1):(1'h0)]) ^~ $signed($unsigned(reg145)))));
            end
          else
            begin
              reg152 <= wire130;
              reg153 <= reg137[(4'he):(4'h8)];
              reg154 <= {wire133,
                  (~((&$unsigned(wire148)) ?
                      (&(reg136 << reg150)) : reg136[(1'h1):(1'h0)]))};
              reg155 <= $unsigned(($signed((wire134[(1'h0):(1'h0)] ^~ $signed(reg151))) != $signed(((reg153 || wire130) < (|reg152)))));
              reg156 <= wire130[(3'h5):(2'h2)];
            end
        end
      else
        begin
          if ($unsigned(reg156[(2'h2):(2'h2)]))
            begin
              reg152 <= reg154;
            end
          else
            begin
              reg152 <= (^~(~&{reg153[(3'h4):(2'h3)]}));
              reg153 <= (reg146 ?
                  $signed(($unsigned($signed(wire133)) ?
                      $signed((~|reg146)) : (~(wire149 ?
                          reg145 : (8'ha6))))) : (8'ha1));
            end
          reg154 <= (&wire130[(4'hb):(4'h9)]);
        end
      if (($unsigned(reg154) ^~ ((!$unsigned((8'hba))) && reg141)))
        begin
          reg157 <= ((8'ha7) ? reg147 : wire138);
          if (reg137)
            begin
              reg158 <= ((reg143 <= $signed(reg153)) ?
                  ($signed(reg140[(4'h8):(2'h2)]) ?
                      (((wire133 << reg155) >= reg144) ?
                          $unsigned((reg154 & reg147)) : $unsigned((wire133 ?
                              reg157 : (8'hb5)))) : wire134[(1'h1):(1'h1)]) : $signed((($signed(reg141) < (~&reg157)) ?
                      $unsigned(wire132[(3'h4):(2'h2)]) : reg145)));
            end
          else
            begin
              reg158 <= $signed({{((~reg157) >>> wire133[(4'ha):(2'h2)])}});
            end
        end
      else
        begin
          reg157 <= ($unsigned(((+$signed((8'ha2))) ?
                  ((reg136 ? reg136 : reg152) ?
                      (reg157 ?
                          wire129 : wire148) : $signed(reg139)) : ((~&reg158) ^ (reg140 << reg141)))) ?
              (^~$unsigned((8'hb2))) : ($unsigned($unsigned({(8'ha5),
                      (8'h9e)})) ?
                  (8'hbc) : (!reg144[(3'h5):(2'h2)])));
          reg158 <= {((((reg139 >>> reg150) > (wire149 <<< wire130)) ?
                      $unsigned($signed(wire138)) : (-(wire135 <= (8'hae)))) ?
                  reg140[(4'hb):(4'h8)] : $signed(reg147)),
              (&reg158)};
          if (reg136)
            begin
              reg159 <= reg155[(3'h6):(3'h4)];
              reg160 <= ((((~|reg150[(3'h5):(2'h3)]) ?
                  $unsigned(wire129[(3'h6):(2'h2)]) : $unsigned(((8'ha1) || (8'h9f)))) ^~ {wire149[(3'h4):(1'h1)]}) || reg146[(4'ha):(2'h2)]);
            end
          else
            begin
              reg159 <= (~^{reg154[(3'h6):(3'h4)],
                  $unsigned({reg143[(2'h3):(1'h1)]})});
              reg160 <= reg147;
              reg161 <= reg146[(4'he):(4'hb)];
            end
        end
      reg162 <= (8'hab);
    end
  assign wire163 = ($signed(reg159[(1'h1):(1'h0)]) ?
                       (!$signed(wire131)) : reg137);
  assign wire164 = {reg160, wire148[(4'h8):(2'h3)]};
  assign wire165 = wire133;
  assign wire166 = (8'h9f);
  assign wire167 = $unsigned(wire149);
  assign wire168 = $unsigned($signed((($unsigned(wire164) >= (reg161 ?
                           reg150 : reg150)) ?
                       reg157 : $signed((+wire129)))));
endmodule