module top  (y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h233):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire0;
  input wire signed [(4'hf):(1'h0)] wire1;
  input wire signed [(5'h15):(1'h0)] wire2;
  input wire signed [(4'h9):(1'h0)] wire3;
  input wire [(5'h10):(1'h0)] wire4;
  reg [(5'h12):(1'h0)] reg414 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire412;
  wire [(4'he):(1'h0)] wire210;
  wire [(5'h12):(1'h0)] wire209;
  wire [(4'hc):(1'h0)] wire208;
  wire [(5'h15):(1'h0)] wire207;
  reg signed [(5'h11):(1'h0)] reg206 = (1'h0);
  reg [(5'h13):(1'h0)] reg205 = (1'h0);
  reg [(5'h14):(1'h0)] reg204 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg203 = (1'h0);
  reg [(5'h15):(1'h0)] reg202 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg201 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar200 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire199;
  reg [(5'h13):(1'h0)] reg198 = (1'h0);
  reg [(3'h4):(1'h0)] reg197 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar196 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg195 = (1'h0);
  wire [(5'h11):(1'h0)] wire194;
  wire [(5'h13):(1'h0)] wire193;
  reg [(5'h11):(1'h0)] reg192 = (1'h0);
  reg [(4'h8):(1'h0)] reg191 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg190 = (1'h0);
  reg [(3'h4):(1'h0)] reg189 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg188 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg187 = (1'h0);
  reg [(4'hc):(1'h0)] reg186 = (1'h0);
  reg [(5'h11):(1'h0)] forvar185 = (1'h0);
  reg [(3'h4):(1'h0)] reg184 = (1'h0);
  reg [(3'h6):(1'h0)] forvar183 = (1'h0);
  reg [(2'h2):(1'h0)] reg182 = (1'h0);
  reg [(4'he):(1'h0)] reg181 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire180;
  wire [(4'ha):(1'h0)] wire179;
  reg [(4'h9):(1'h0)] reg178 = (1'h0);
  reg [(4'hf):(1'h0)] reg177 = (1'h0);
  reg [(4'hf):(1'h0)] reg176 = (1'h0);
  reg [(3'h4):(1'h0)] reg175 = (1'h0);
  reg [(3'h4):(1'h0)] forvar174 = (1'h0);
  reg [(5'h15):(1'h0)] reg173 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg172 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg171 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg170 = (1'h0);
  wire [(4'ha):(1'h0)] wire169;
  wire signed [(4'hb):(1'h0)] wire5;
  wire signed [(3'h6):(1'h0)] wire167;
  assign y = {reg414,
                 wire412,
                 wire210,
                 wire209,
                 wire208,
                 wire207,
                 reg206,
                 reg205,
                 reg204,
                 reg203,
                 reg202,
                 reg201,
                 forvar200,
                 wire199,
                 reg198,
                 reg197,
                 forvar196,
                 reg195,
                 wire194,
                 wire193,
                 reg192,
                 reg191,
                 reg190,
                 reg189,
                 reg188,
                 reg187,
                 reg186,
                 forvar185,
                 reg184,
                 forvar183,
                 reg182,
                 reg181,
                 wire180,
                 wire179,
                 reg178,
                 reg177,
                 reg176,
                 reg175,
                 forvar174,
                 reg173,
                 reg172,
                 reg171,
                 reg170,
                 wire169,
                 wire5,
                 wire167,
                 (1'h0)};
  assign wire5 = wire1;
  module6 modinst168 (.wire8(wire4), .wire10(wire1), .wire7(wire0), .wire11(wire3), .y(wire167), .wire9(wire5), .clk(clk));
  assign wire169 = wire167;
  always
    @(posedge clk) begin
      reg170 = ((wire3 || {wire1, wire1}) ?
          $unsigned(wire0) : wire169[(3'h6):(1'h0)]);
      reg171 <= $unsigned((-wire4));
      reg172 <= (wire4[(4'hf):(4'hf)] > $signed({{wire4[(3'h4):(2'h3)]}}));
    end
  always
    @(posedge clk) begin
      reg173 <= ($unsigned($signed($signed((wire2 ? wire169 : (8'hac))))) ?
          $unsigned(((|(!(8'haa))) ?
              reg171 : $unsigned($signed(wire5)))) : (~$signed({(^wire2),
              $unsigned(wire3)})));
      reg177 <= $signed(({(8'hbe), wire4[(3'h4):(3'h4)]} ?
          (+wire1) : ($signed((+wire4)) >> {(wire1 ? forvar174 : forvar174),
              ((8'hb7) * reg176)})));
      reg178 <= {($signed(forvar174[(1'h0):(1'h0)]) ?
              ((&(~&(8'hb7))) >> $unsigned((reg171 ^ reg175))) : wire2[(4'hd):(1'h0)])};
    end
  assign wire179 = ((~|wire167[(3'h5):(2'h3)]) ? reg172 : $unsigned(wire169));
  assign wire180 = ((((~|(reg175 <<< wire1)) | $signed((reg178 >= reg171))) ?
                           ($signed($unsigned(reg176)) < reg172) : ($signed((7'h43)) ~^ wire179[(3'h5):(2'h3)])) ?
                       (wire179[(3'h4):(2'h2)] ?
                           reg170[(3'h5):(1'h0)] : wire179) : forvar174[(2'h2):(2'h2)]);
  always
    @(posedge clk) begin
      reg181 <= (~forvar174);
      reg182 = ($unsigned((reg175 ?
              $unsigned((~&wire169)) : $unsigned($signed((8'hb9))))) ?
          (~|{reg177, (|wire167)}) : $unsigned(wire4));
      for (forvar183 = (1'h0); (forvar183 < (1'h1)); forvar183 = (forvar183 + (1'h1)))
        begin
          reg184 = $unsigned(wire167[(1'h0):(1'h0)]);
          for (forvar185 = (1'h0); (forvar185 < (2'h2)); forvar185 = (forvar185 + (1'h1)))
            begin
              reg186 <= reg176;
              reg187 = (|$unsigned((~(^((8'hb2) ? wire4 : wire0)))));
              reg188 <= (wire0 ?
                  $signed(wire179) : (($unsigned((wire5 ? reg170 : reg172)) ?
                      (~reg173[(1'h1):(1'h0)]) : (|(~|wire180))) * ({(&(8'hb3)),
                      (reg172 < wire169)} || ($signed(reg170) == $signed(wire167)))));
              reg189 <= ($signed(((~^((7'h44) ? (8'hbe) : forvar183)) ?
                  wire169[(3'h7):(1'h0)] : (-(reg181 <<< reg178)))) | forvar183[(1'h0):(1'h0)]);
              reg190 <= $unsigned(wire3);
            end
          reg191 <= (+($unsigned(reg187) << ((reg187[(3'h6):(3'h5)] ?
              wire180[(4'ha):(2'h2)] : {wire3}) || (~^reg173))));
        end
      reg192 <= $signed((8'hab));
    end
  assign wire193 = wire180[(4'ha):(1'h1)];
  assign wire194 = {(&wire3[(3'h7):(3'h4)]),
                       ($unsigned(({reg182,
                           reg189} ^~ {(7'h44)})) <<< $signed({(reg170 - (8'hae)),
                           $unsigned(reg177)}))};
  always
    @(posedge clk) begin
      reg195 <= reg188[(2'h3):(2'h3)];
      for (forvar196 = (1'h0); (forvar196 < (2'h3)); forvar196 = (forvar196 + (1'h1)))
        begin
          reg197 <= reg182;
          reg198 <= reg187;
        end
    end
  assign wire199 = (8'hac);
  always
    @(posedge clk) begin
      for (forvar200 = (1'h0); (forvar200 < (2'h3)); forvar200 = (forvar200 + (1'h1)))
        begin
          reg201 = reg186[(2'h2):(2'h2)];
          reg202 <= {(8'hb4), reg173};
          reg203 <= forvar183[(3'h6):(3'h4)];
          reg204 = $signed((((~&$signed((8'h9c))) ?
              (8'had) : ((wire3 && wire180) - (~^wire0))) && $unsigned(reg172[(1'h1):(1'h1)])));
          reg205 = (forvar200[(4'hc):(1'h1)] ?
              ((8'hbc) <<< {wire4}) : (($signed((~|wire4)) - wire3) ?
                  $unsigned(reg190[(4'hb):(3'h4)]) : $signed(wire194)));
        end
      reg206 = $signed(($unsigned((reg181 | reg175)) ?
          (^~$signed(reg190)) : $unsigned({$unsigned(forvar185),
              (&forvar196)})));
    end
  assign wire207 = forvar174[(2'h2):(1'h0)];
  assign wire208 = (({wire180} ?
                           wire169[(4'ha):(4'h9)] : ((((8'had) >> reg206) ?
                               (7'h42) : wire2[(5'h15):(3'h4)]) && $unsigned($signed(wire179)))) ?
                       ((((8'h9c) ? reg177 : (reg203 ? wire180 : (8'hbf))) ?
                               ({forvar185} ?
                                   (8'hbf) : (!reg188)) : $unsigned(wire169[(3'h7):(2'h3)])) ?
                           $unsigned($signed({reg205})) : (~^(reg191 > (~&reg173)))) : (8'ha9));
  assign wire209 = reg175[(1'h0):(1'h0)];
  assign wire210 = $signed($unsigned($unsigned({(|(8'h9e)),
                       $unsigned((8'hb0))})));
  module211 modinst413 (.wire214(reg173), .clk(clk), .y(wire412), .wire215(reg195), .wire212(forvar196), .wire213(wire180));
  always
    @(posedge clk) begin
      reg414 <= $unsigned($unsigned((~&((forvar174 ?
          wire199 : forvar200) && {reg206, wire209}))));
    end
endmodule

module module211
#( parameter param411 = (^~((((!(8'hba)) < ((8'ha7) * (8'hae))) ? (((8'hb2) - (8'hbc)) ? ((8'hbb) ? (8'ha3) : (8'had)) : ((7'h42) ? (8'hb7) : (8'h9c))) : (~|((8'hb1) ? (8'h9c) : (8'hb3)))) ? {(((8'ha3) && (8'hb3)) ~^ (&(8'ha0)))} : ((!((8'hba) & (8'h9f))) ? ({(8'hbe), (8'hb2)} ? ((8'ha6) + (8'hb9)) : (~(8'hbd))) : (-((8'hb7) >>> (8'hba)))))) )
(y, clk, wire212, wire213, wire214, wire215);
  output wire [(32'h148):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire212;
  input wire signed [(4'h9):(1'h0)] wire213;
  input wire signed [(5'h15):(1'h0)] wire214;
  input wire [(3'h7):(1'h0)] wire215;
  wire [(3'h5):(1'h0)] wire410;
  wire [(2'h3):(1'h0)] wire408;
  reg [(2'h2):(1'h0)] reg274 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg273 = (1'h0);
  reg [(4'hc):(1'h0)] reg272 = (1'h0);
  reg [(4'hc):(1'h0)] reg271 = (1'h0);
  reg [(5'h12):(1'h0)] reg270 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg269 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg268 = (1'h0);
  reg [(3'h4):(1'h0)] forvar267 = (1'h0);
  wire [(4'hc):(1'h0)] wire266;
  reg signed [(3'h5):(1'h0)] reg265 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg264 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg263 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire262;
  wire signed [(5'h12):(1'h0)] wire261;
  reg [(5'h10):(1'h0)] reg216 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg217 = (1'h0);
  reg [(4'hf):(1'h0)] reg218 = (1'h0);
  reg [(2'h2):(1'h0)] reg219 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg220 = (1'h0);
  reg [(3'h4):(1'h0)] reg221 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg222 = (1'h0);
  reg [(3'h7):(1'h0)] forvar223 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg224 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar225 = (1'h0);
  reg [(4'h9):(1'h0)] reg226 = (1'h0);
  reg [(4'he):(1'h0)] reg227 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg228 = (1'h0);
  reg [(4'hc):(1'h0)] reg229 = (1'h0);
  reg [(4'hf):(1'h0)] reg230 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire259;
  assign y = {wire410,
                 wire408,
                 reg274,
                 reg273,
                 reg272,
                 reg271,
                 reg270,
                 reg269,
                 reg268,
                 forvar267,
                 wire266,
                 reg265,
                 reg264,
                 reg263,
                 wire262,
                 wire261,
                 reg216,
                 reg217,
                 reg218,
                 reg219,
                 reg220,
                 reg221,
                 reg222,
                 forvar223,
                 reg224,
                 forvar225,
                 reg226,
                 reg227,
                 reg228,
                 reg229,
                 reg230,
                 wire259,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg216 <= ($unsigned((^{$unsigned((8'hb9))})) ?
          (^(wire215[(3'h4):(2'h2)] | wire214)) : $unsigned($unsigned(wire212)));
      reg217 <= reg216;
      reg218 <= reg217[(3'h6):(2'h3)];
    end
  always
    @(posedge clk) begin
      reg219 <= $signed($signed(($signed(wire213[(2'h2):(1'h0)]) & $signed($unsigned(reg218)))));
      reg220 <= $signed((reg217 * (($unsigned(wire214) ?
              {wire215} : (|reg219)) ?
          $unsigned((reg217 * reg216)) : {(wire214 ? wire215 : reg216)})));
      reg221 <= (|wire212);
      reg222 <= reg217[(3'h7):(3'h5)];
      for (forvar223 = (1'h0); (forvar223 < (2'h3)); forvar223 = (forvar223 + (1'h1)))
        begin
          reg224 <= wire215[(1'h0):(1'h0)];
          for (forvar225 = (1'h0); (forvar225 < (1'h1)); forvar225 = (forvar225 + (1'h1)))
            begin
              reg226 <= (reg219 & ($unsigned($unsigned(((8'h9c) ?
                  reg218 : forvar223))) * {($unsigned(reg221) ?
                      $signed(wire213) : $signed((7'h41)))}));
              reg227 = reg216;
              reg228 = reg220;
              reg229 <= ($unsigned((reg217 && ((reg220 + wire214) ?
                      (+reg228) : (reg222 <<< reg216)))) ?
                  (~&reg227[(2'h3):(2'h2)]) : $signed(forvar223[(3'h6):(1'h0)]));
              reg230 <= (forvar223 ^ (!((+{wire215}) - $signed({wire215,
                  (8'ha3)}))));
            end
        end
    end
  module231 modinst260 (.wire233(reg218), .y(wire259), .wire232(reg226), .wire235(reg221), .wire234(reg230), .clk(clk), .wire236(reg227));
  assign wire261 = (forvar223 ?
                       (wire213 ?
                           {$unsigned((wire215 ^~ (7'h44)))} : $unsigned($signed(wire259))) : ((reg219 ^ $signed(((8'ha5) ^~ reg222))) <= (-wire214[(4'h8):(3'h5)])));
  assign wire262 = reg221;
  always
    @(posedge clk) begin
      reg263 <= (8'ha3);
    end
  always
    @(posedge clk) begin
      reg264 = $unsigned(reg224);
    end
  always
    @(posedge clk) begin
      reg265 <= ($unsigned(forvar225) ?
          (8'ha3) : ($unsigned($signed(reg229)) ?
              wire261[(5'h10):(5'h10)] : $signed($unsigned($signed((8'h9e))))));
    end
  assign wire266 = wire262[(3'h7):(3'h4)];
  always
    @(posedge clk) begin
      for (forvar267 = (1'h0); (forvar267 < (2'h2)); forvar267 = (forvar267 + (1'h1)))
        begin
          reg268 <= $unsigned(reg264[(1'h0):(1'h0)]);
          reg269 = (8'hbd);
          reg270 <= $unsigned($signed($unsigned(wire262)));
          reg271 = ((((~|$unsigned(reg217)) && $signed(reg218[(4'hc):(3'h4)])) ?
              (~^wire212) : (((reg268 ? wire266 : reg229) == $signed(reg229)) ?
                  ({reg229} ?
                      (wire212 ^ reg217) : (forvar267 ?
                          reg221 : reg217)) : reg224[(3'h6):(1'h1)])) ^ {reg218[(3'h6):(1'h1)]});
        end
      reg272 <= (($signed(($signed((8'hb5)) ?
              {wire212, (8'hb0)} : $signed(reg263))) * wire261) ?
          ($unsigned(wire261) + $unsigned(forvar267)) : ((~^$unsigned((forvar223 != forvar225))) ?
              ((reg270 != (^~reg218)) ?
                  $unsigned($unsigned(forvar267)) : reg265) : (8'ha1)));
      reg273 = $unsigned($signed(wire262));
      reg274 <= (reg217[(4'hd):(3'h6)] ?
          ((reg226[(2'h2):(1'h1)] * ((wire261 ? (8'hb6) : reg272) ?
                  (wire262 ^ wire215) : (8'hbf))) ?
              $unsigned(reg271[(4'hb):(3'h6)]) : wire266) : wire215);
    end
  module275 modinst409 (.wire279(reg226), .wire278(wire213), .wire276(wire214), .y(wire408), .clk(clk), .wire277(wire261));
  assign wire410 = reg224;
endmodule

module module6
#( parameter param166 = (({{((8'hb7) - (8'ha1))}, (((8'hb8) ? (8'h9e) : (8'hb5)) ? (^(8'hb4)) : (~&(8'h9f)))} ^~ {(^~((8'h9f) ? (8'ha0) : (8'ha7)))}) ? (8'h9c) : ((8'hb8) == {(((8'ha1) | (8'hae)) ? (~&(8'haa)) : (-(8'ha5)))})) )
(y, clk, wire7, wire8, wire9, wire10, wire11);
  output wire [(32'ha5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire7;
  input wire signed [(4'hc):(1'h0)] wire8;
  input wire [(4'hb):(1'h0)] wire9;
  input wire signed [(4'h8):(1'h0)] wire10;
  input wire signed [(4'h9):(1'h0)] wire11;
  reg [(4'hb):(1'h0)] reg165 = (1'h0);
  reg [(2'h2):(1'h0)] reg164 = (1'h0);
  reg [(5'h15):(1'h0)] reg163 = (1'h0);
  wire [(4'h9):(1'h0)] wire162;
  reg signed [(5'h15):(1'h0)] reg161 = (1'h0);
  wire [(5'h11):(1'h0)] wire12;
  wire signed [(4'hc):(1'h0)] wire13;
  reg [(3'h4):(1'h0)] reg14 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg15 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg16 = (1'h0);
  reg [(4'hf):(1'h0)] reg17 = (1'h0);
  reg [(4'hc):(1'h0)] reg18 = (1'h0);
  wire [(4'hb):(1'h0)] wire159;
  assign y = {reg165,
                 reg164,
                 reg163,
                 wire162,
                 reg161,
                 wire12,
                 wire13,
                 reg14,
                 reg15,
                 reg16,
                 reg17,
                 reg18,
                 wire159,
                 (1'h0)};
  assign wire12 = ((({(wire11 * wire9), wire9[(4'h9):(2'h3)]} ?
                              wire8[(2'h2):(1'h0)] : wire7) ?
                          $signed(wire9) : $signed((|(~|wire8)))) ?
                      $unsigned((wire7[(3'h5):(3'h5)] + $signed((wire11 + wire7)))) : wire11[(2'h2):(1'h1)]);
  assign wire13 = $signed(wire8[(2'h2):(1'h0)]);
  always
    @(posedge clk) begin
      reg14 <= {$unsigned($unsigned(wire9[(3'h7):(1'h1)]))};
      reg15 <= ({(~|((reg14 ? (8'h9f) : wire7) ^ $signed(reg14))),
          {$unsigned((wire13 ?
                  wire12 : wire9))}} ^ $unsigned({wire13[(4'ha):(1'h0)],
          ($unsigned(wire11) ? (&(8'hb7)) : wire10)}));
      reg16 <= $signed(wire8);
      reg17 = ($signed(wire12[(4'he):(4'h8)]) | wire11);
      reg18 <= $signed((wire11[(3'h7):(1'h0)] ? (+wire13) : wire7));
    end
  module19 modinst160 (wire159, clk, reg16, wire7, wire10, wire9, reg15);
  always
    @(posedge clk) begin
      reg161 <= $unsigned((reg18 ?
          reg15[(3'h4):(1'h1)] : $signed(((wire11 ? (8'hb9) : wire8) ?
              ((8'hbe) | wire11) : $signed(wire9)))));
    end
  assign wire162 = wire9;
  always
    @(posedge clk) begin
      reg163 = wire10[(3'h4):(1'h1)];
    end
  always
    @(posedge clk) begin
      reg164 <= (($unsigned($signed((reg16 ? (8'haa) : (8'hb5)))) ?
              {$signed((~&wire8)), $unsigned($signed(wire12))} : (8'hbe)) ?
          {($unsigned((reg17 == (8'ha5))) ~^ (&(wire7 ? wire7 : reg18))),
              (wire9 ?
                  (&(wire13 + wire8)) : (~(reg14 >> reg18)))} : $unsigned((((7'h40) == (wire159 ?
              wire10 : reg161)) ^ reg15[(4'h9):(2'h3)])));
      reg165 <= ({reg163} ?
          ((!reg16) ^ $unsigned(wire162[(3'h6):(1'h1)])) : wire10);
    end
endmodule

module module19
#( parameter param158 = (({((~|(8'hbf)) ^ ((8'hbc) || (8'hb6)))} ? ({{(8'hbd)}, (8'hb9)} ? {((8'hab) ? (8'hbb) : (8'hb9)), ((8'hb5) & (8'hbe))} : ({(8'haf), (8'hb8)} ? ((8'ha8) * (7'h44)) : (!(8'hba)))) : (~(|(+(8'hbf))))) > {((~|{(8'ha7), (8'hb6)}) ^~ (((8'hab) ? (7'h43) : (8'hbe)) && ((7'h42) ^~ (8'hbe)))), ((~&{(8'ha0), (8'ha4)}) ? {{(8'h9f), (8'hbf)}, (!(7'h41))} : (((8'hb2) == (8'haf)) - ((8'hb8) ? (8'hbf) : (8'hb1))))}) )
(y, clk, wire24, wire23, wire22, wire21, wire20);
  output wire [(32'h1b0):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire24;
  input wire [(4'he):(1'h0)] wire23;
  input wire signed [(4'h8):(1'h0)] wire22;
  input wire signed [(3'h5):(1'h0)] wire21;
  input wire signed [(3'h7):(1'h0)] wire20;
  wire [(5'h13):(1'h0)] wire157;
  wire [(4'hd):(1'h0)] wire78;
  wire [(4'hd):(1'h0)] wire38;
  reg [(5'h11):(1'h0)] reg37 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg36 = (1'h0);
  reg [(4'hf):(1'h0)] reg35 = (1'h0);
  reg [(4'hf):(1'h0)] reg34 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg33 = (1'h0);
  reg [(4'ha):(1'h0)] forvar32 = (1'h0);
  wire [(3'h7):(1'h0)] wire31;
  wire signed [(4'hb):(1'h0)] wire30;
  wire [(4'hf):(1'h0)] wire29;
  wire [(4'hd):(1'h0)] wire28;
  wire signed [(5'h14):(1'h0)] wire27;
  reg signed [(4'hb):(1'h0)] reg26 = (1'h0);
  reg [(5'h12):(1'h0)] reg25 = (1'h0);
  wire [(3'h5):(1'h0)] wire80;
  wire [(3'h6):(1'h0)] wire81;
  wire [(4'hd):(1'h0)] wire82;
  reg [(4'h8):(1'h0)] forvar83 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar84 = (1'h0);
  reg [(3'h6):(1'h0)] reg85 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg86 = (1'h0);
  reg [(4'hb):(1'h0)] reg87 = (1'h0);
  reg [(4'he):(1'h0)] reg88 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg89 = (1'h0);
  reg [(4'hd):(1'h0)] reg90 = (1'h0);
  reg [(4'hc):(1'h0)] reg91 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg92 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg93 = (1'h0);
  wire [(5'h13):(1'h0)] wire94;
  reg [(3'h7):(1'h0)] reg95 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg96 = (1'h0);
  wire [(4'hd):(1'h0)] wire155;
  assign y = {wire157,
                 wire78,
                 wire38,
                 reg37,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 forvar32,
                 wire31,
                 wire30,
                 wire29,
                 wire28,
                 wire27,
                 reg26,
                 reg25,
                 wire80,
                 wire81,
                 wire82,
                 forvar83,
                 forvar84,
                 reg85,
                 reg86,
                 reg87,
                 reg88,
                 reg89,
                 reg90,
                 reg91,
                 reg92,
                 reg93,
                 wire94,
                 reg95,
                 reg96,
                 wire155,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg25 <= $signed($unsigned((($signed((8'hb2)) ?
          $unsigned(wire24) : $signed(wire20)) << ($unsigned(wire23) || wire24[(4'hb):(2'h3)]))));
      reg26 = (wire21[(2'h2):(1'h0)] ?
          ($signed(((reg25 ?
              wire20 : wire24) * wire20[(2'h2):(1'h1)])) && (((wire21 >>> wire20) * (wire22 <<< wire20)) ?
              wire23 : (~^{(8'ha0), (8'hbb)}))) : wire23[(3'h4):(2'h2)]);
    end
  assign wire27 = (reg25 ?
                      (wire23[(2'h2):(1'h1)] - reg25[(3'h4):(3'h4)]) : wire21[(1'h0):(1'h0)]);
  assign wire28 = {$unsigned(({wire21} ?
                          ((8'hb0) * wire24[(5'h10):(2'h3)]) : wire20))};
  assign wire29 = $unsigned(((|(!wire21)) ?
                      wire22 : (($unsigned(wire24) ?
                          wire22 : (wire22 < wire21)) && $signed((~|wire22)))));
  assign wire30 = wire24[(4'hc):(2'h3)];
  assign wire31 = ($signed({wire23}) ?
                      (~&wire28[(3'h4):(1'h1)]) : (~(&((8'hb5) >>> (^wire20)))));
  always
    @(posedge clk) begin
      for (forvar32 = (1'h0); (forvar32 < (1'h1)); forvar32 = (forvar32 + (1'h1)))
        begin
          reg33 <= ($signed(wire29[(3'h7):(2'h2)]) ?
              (&((&{wire22, wire27}) ?
                  $signed({(8'h9d)}) : $unsigned((wire23 <<< reg25)))) : (~&(&wire28)));
          reg34 <= (~^(wire27[(4'he):(4'he)] + forvar32));
        end
      reg35 = wire28[(4'h8):(4'h8)];
      reg36 = (7'h41);
      reg37 <= (reg35 ?
          ($unsigned(((reg34 > (8'hb0)) - (wire24 ^ reg25))) ^ (~^forvar32)) : $unsigned($signed(reg36)));
    end
  assign wire38 = ((&{$unsigned(((7'h42) != reg26))}) ?
                      (((8'ha8) ?
                          reg35[(4'hb):(4'h8)] : ($unsigned(forvar32) ?
                              (!reg35) : reg37)) - $unsigned(($signed(wire31) <<< wire22[(3'h4):(1'h1)]))) : wire27);
  module39 modinst79 (wire78, clk, wire29, reg26, reg25, reg36, reg34);
  assign wire80 = ((~($signed($unsigned(wire22)) ?
                          $signed((forvar32 ?
                              wire23 : forvar32)) : ((wire21 <= reg35) || reg25[(1'h1):(1'h1)]))) ?
                      $signed($signed((wire28[(2'h2):(1'h0)] >>> (^~reg26)))) : $unsigned((reg36[(3'h5):(3'h5)] <<< $unsigned(wire27[(3'h7):(1'h0)]))));
  assign wire81 = (~(reg36[(4'h8):(3'h4)] >= (wire80 ?
                      (8'hb9) : $signed($unsigned(reg36)))));
  assign wire82 = ($signed((((+wire23) ?
                          wire80[(1'h0):(1'h0)] : (wire24 | reg35)) ?
                      $unsigned((~|wire38)) : reg33[(1'h0):(1'h0)])) <<< {((reg25[(4'he):(4'h9)] ?
                              (wire21 || reg36) : {wire23}) ?
                          {(wire24 <<< wire29),
                              {wire30}} : (reg35 == (wire28 > reg35))),
                      {(forvar32[(3'h6):(2'h2)] <= $signed(wire31))}});
  always
    @(posedge clk) begin
      for (forvar83 = (1'h0); (forvar83 < (2'h3)); forvar83 = (forvar83 + (1'h1)))
        begin
          for (forvar84 = (1'h0); (forvar84 < (1'h1)); forvar84 = (forvar84 + (1'h1)))
            begin
              reg85 = wire82[(4'hd):(4'ha)];
              reg86 <= $unsigned((8'hb1));
              reg87 <= $signed({$signed(reg35[(4'hc):(1'h0)]), wire38});
              reg88 <= (8'ha1);
            end
          reg89 <= $unsigned((^$unsigned(wire82[(4'hd):(4'ha)])));
          reg90 <= (^$unsigned((~|($signed(wire82) ?
              (wire82 ? reg26 : reg35) : ((8'h9d) ? wire80 : reg36)))));
        end
      reg91 <= (8'hbc);
      reg92 <= ($signed((wire23 ?
              {$signed(wire31)} : ($unsigned(reg36) * (wire82 ?
                  forvar83 : wire30)))) ?
          (reg35 ^ $unsigned(((wire78 ?
              wire81 : reg90) ^ $unsigned(wire78)))) : wire20);
      reg93 = forvar84[(4'ha):(1'h0)];
    end
  assign wire94 = (((({reg91,
                              wire20} << {forvar83}) <= (reg92[(4'h9):(1'h0)] == $signed(reg37))) ?
                          $unsigned({reg86[(3'h6):(2'h2)]}) : reg35[(3'h5):(2'h3)]) ?
                      ({(&{reg89})} >> ($unsigned(wire30) ?
                          $unsigned(wire27) : {(wire78 ? wire28 : wire81),
                              (reg36 ?
                                  reg91 : wire29)})) : ($unsigned(((reg34 >= reg36) ?
                          wire78[(4'hb):(3'h7)] : (wire23 ?
                              (8'h9d) : forvar32))) ^~ (^{$signed(wire31)})));
  always
    @(posedge clk) begin
      reg95 <= $signed(wire23[(3'h5):(2'h2)]);
      reg96 <= (((($unsigned(reg33) ?
              (reg85 ^ wire27) : (wire78 ?
                  reg35 : reg35)) != wire78[(2'h3):(2'h2)]) ?
          ($unsigned(wire24[(1'h0):(1'h0)]) >= wire27) : {wire31,
              reg89[(2'h2):(2'h2)]}) >> (~^$unsigned($signed(wire22[(3'h5):(3'h5)]))));
    end
  module97 modinst156 (wire155, clk, wire94, wire21, reg35, wire38, wire24);
  assign wire157 = {$unsigned($unsigned(wire81)), (8'h9e)};
endmodule

module module97  (y, clk, wire102, wire101, wire100, wire99, wire98);
  output wire [(32'h252):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h13):(1'h0)] wire102;
  input wire signed [(2'h3):(1'h0)] wire101;
  input wire [(4'ha):(1'h0)] wire100;
  input wire signed [(4'hd):(1'h0)] wire99;
  input wire [(5'h14):(1'h0)] wire98;
  reg signed [(4'hc):(1'h0)] reg154 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg153 = (1'h0);
  reg [(4'h8):(1'h0)] reg152 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg151 = (1'h0);
  wire [(3'h6):(1'h0)] wire150;
  reg [(2'h2):(1'h0)] reg149 = (1'h0);
  reg [(4'hd):(1'h0)] reg148 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire147;
  wire [(4'hf):(1'h0)] wire146;
  wire signed [(3'h6):(1'h0)] wire145;
  reg [(2'h2):(1'h0)] reg144 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg143 = (1'h0);
  reg [(5'h11):(1'h0)] reg142 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg141 = (1'h0);
  reg [(4'h8):(1'h0)] reg140 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg139 = (1'h0);
  reg [(3'h7):(1'h0)] reg138 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg137 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg136 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar135 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg134 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire133;
  reg [(3'h5):(1'h0)] reg132 = (1'h0);
  reg [(4'he):(1'h0)] reg131 = (1'h0);
  reg [(5'h11):(1'h0)] reg130 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg129 = (1'h0);
  reg [(5'h10):(1'h0)] reg128 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar127 = (1'h0);
  reg signed [(4'he):(1'h0)] reg126 = (1'h0);
  reg [(5'h14):(1'h0)] reg125 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg124 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg123 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg122 = (1'h0);
  reg [(5'h10):(1'h0)] reg121 = (1'h0);
  reg [(3'h5):(1'h0)] reg120 = (1'h0);
  reg [(4'hd):(1'h0)] reg119 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg118 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg117 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg116 = (1'h0);
  reg [(4'hb):(1'h0)] reg115 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg114 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg113 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg112 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg111 = (1'h0);
  reg [(5'h10):(1'h0)] forvar110 = (1'h0);
  reg [(4'h9):(1'h0)] reg109 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg108 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg107 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg106 = (1'h0);
  reg [(5'h14):(1'h0)] forvar105 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg104 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg103 = (1'h0);
  assign y = {reg154,
                 reg153,
                 reg152,
                 reg151,
                 wire150,
                 reg149,
                 reg148,
                 wire147,
                 wire146,
                 wire145,
                 reg144,
                 reg143,
                 reg142,
                 reg141,
                 reg140,
                 reg139,
                 reg138,
                 reg137,
                 reg136,
                 forvar135,
                 reg134,
                 wire133,
                 reg132,
                 reg131,
                 reg130,
                 reg129,
                 reg128,
                 forvar127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 reg117,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 reg112,
                 reg111,
                 forvar110,
                 reg109,
                 reg108,
                 reg107,
                 reg106,
                 forvar105,
                 reg104,
                 reg103,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg103 <= ((wire98[(2'h2):(2'h2)] <= wire99[(4'hd):(4'h9)]) ?
          $signed({($signed(wire99) * wire102[(1'h1):(1'h0)]),
              $signed((~wire100))}) : ((|(8'hba)) ?
              (~&$unsigned((wire102 ? wire102 : wire100))) : (&((^wire98) ?
                  (wire100 || wire98) : wire102[(5'h11):(4'h9)]))));
      reg104 <= (^{$unsigned($signed((+(8'ha2)))), wire102});
      for (forvar105 = (1'h0); (forvar105 < (1'h1)); forvar105 = (forvar105 + (1'h1)))
        begin
          reg106 <= $unsigned(wire100[(3'h6):(3'h6)]);
          reg107 <= $unsigned(wire98[(1'h0):(1'h0)]);
          reg108 <= $signed((wire99 != (reg106[(3'h4):(2'h2)] > reg106[(2'h3):(2'h3)])));
          reg109 <= (+{{$unsigned(wire100[(4'h8):(3'h4)])}, reg107});
          for (forvar110 = (1'h0); (forvar110 < (3'h4)); forvar110 = (forvar110 + (1'h1)))
            begin
              reg111 <= ($signed((wire102[(3'h4):(2'h2)] < $signed($unsigned((7'h40))))) ?
                  reg106 : (-({$unsigned(forvar105),
                      wire100} || reg104[(1'h0):(1'h0)])));
              reg112 <= reg107[(4'hb):(4'hb)];
              reg113 <= (|((-((&wire100) | (reg108 ?
                  reg103 : reg106))) | $signed(((reg108 ~^ (8'hb8)) ?
                  (forvar105 ? reg108 : reg109) : $unsigned(wire101)))));
            end
        end
    end
  always
    @(posedge clk) begin
      reg114 <= reg103;
      reg115 <= $signed(({(|(^reg113))} ?
          (reg112[(2'h2):(1'h0)] + {(reg104 && reg108),
              (wire102 >>> reg109)}) : reg111));
    end
  always
    @(posedge clk) begin
      reg116 <= $signed($signed(((-$signed(reg115)) <<< {{reg108}})));
    end
  always
    @(posedge clk) begin
      reg117 <= {$signed($signed({$signed((8'hbb)), reg115[(4'h8):(1'h1)]}))};
      reg118 = ((reg115 < (((reg116 ?
                  wire99 : wire98) || (forvar110 >>> wire100)) ?
              ((~(7'h44)) == (!forvar110)) : ((reg108 ^ reg106) ?
                  $signed(reg112) : $unsigned(wire102)))) ?
          $unsigned(reg103) : wire99[(3'h6):(3'h5)]);
      reg119 = ({$signed((forvar110[(4'hd):(3'h6)] ? {reg104} : reg106)),
              $signed($unsigned({wire102, reg112}))} ?
          wire102 : $signed($signed(($unsigned(reg103) ^ wire99[(4'h9):(2'h2)]))));
      reg120 = ({$unsigned({$unsigned(reg109), (wire98 | reg106)}),
              reg103[(1'h0):(1'h0)]} ?
          ((~&({reg118, reg118} + (reg113 ? wire100 : reg114))) ?
              $signed((^~(wire102 >= reg106))) : (((forvar110 ~^ reg108) == (^~reg107)) >= {{reg113}})) : (reg119 ?
              $signed($unsigned($unsigned(reg106))) : (~|($signed(reg111) > reg119[(2'h2):(1'h1)]))));
    end
  always
    @(posedge clk) begin
      reg121 <= ((~&(forvar110 ?
              $unsigned(reg113) : ((reg114 == reg120) && $unsigned(forvar110)))) ?
          $signed((8'ha3)) : {$unsigned(({reg115} || reg106))});
    end
  always
    @(posedge clk) begin
      reg122 <= (+(-(-reg116)));
      reg123 <= ($signed(wire102) && reg120[(3'h5):(2'h2)]);
      reg124 <= reg107;
      reg125 <= ((7'h41) | $unsigned(wire98[(3'h6):(2'h2)]));
    end
  always
    @(posedge clk) begin
      reg126 = $signed($signed(({$signed(forvar110), wire102[(4'hc):(4'ha)]} ?
          ($signed(wire99) ?
              (|reg107) : $unsigned(wire100)) : $unsigned((!reg114)))));
      for (forvar127 = (1'h0); (forvar127 < (3'h4)); forvar127 = (forvar127 + (1'h1)))
        begin
          reg128 = $unsigned($unsigned($unsigned($unsigned($unsigned(reg106)))));
          reg129 <= wire98[(3'h7):(3'h5)];
          reg130 <= ({$signed(wire99[(4'h8):(3'h5)]),
                  (~&(~&$signed((8'ha0))))} ?
              $unsigned($unsigned($signed((reg116 ?
                  wire100 : forvar127)))) : reg125);
          reg131 <= ($signed($signed((~forvar110))) < $unsigned((reg125[(2'h2):(1'h1)] ?
              {(~reg124), reg129[(3'h6):(3'h5)]} : reg113[(3'h4):(2'h2)])));
        end
      reg132 = reg103;
    end
  assign wire133 = $signed((8'hb5));
  always
    @(posedge clk) begin
      reg134 <= {$signed($signed({$unsigned((8'ha2)), (reg107 && reg120)})),
          $unsigned(forvar110)};
      for (forvar135 = (1'h0); (forvar135 < (2'h2)); forvar135 = (forvar135 + (1'h1)))
        begin
          reg136 <= reg106[(3'h4):(3'h4)];
          reg137 <= reg129[(4'h9):(1'h1)];
          reg138 <= (reg123 - reg112);
          reg139 = reg119[(4'h9):(4'h8)];
          if ($unsigned(forvar105[(4'hc):(4'hc)]))
            begin
              reg140 <= reg118;
              reg141 <= ($unsigned($unsigned($signed((-(8'hb9))))) ?
                  $unsigned($signed($unsigned($signed(reg120)))) : reg122[(4'hc):(1'h1)]);
              reg142 = (reg132 ? reg131[(4'hd):(3'h5)] : {(8'h9e)});
              reg143 <= (((~&$unsigned(reg119[(1'h1):(1'h1)])) ?
                      (($signed(wire100) ?
                          (-reg137) : (reg106 ?
                              forvar110 : (8'ha4))) || (wire98 ?
                          $signed(wire101) : (+reg115))) : $unsigned(($unsigned(reg132) ?
                          $signed(reg137) : $unsigned(reg109)))) ?
                  reg111[(1'h0):(1'h0)] : $signed(reg104));
              reg144 <= $unsigned((-($unsigned((|reg131)) && {((8'haa) ?
                      reg128 : reg122),
                  ((8'hae) != reg122)})));
            end
          else
            begin
              reg140 = reg141[(1'h0):(1'h0)];
              reg141 <= $unsigned(((-reg142[(4'hd):(4'h8)]) >>> ((~|reg130[(3'h7):(3'h6)]) ?
                  $signed((reg138 ?
                      (7'h40) : reg124)) : (^~(forvar105 ^ reg104)))));
              reg142 <= wire100;
            end
        end
    end
  assign wire145 = reg108;
  assign wire146 = (wire133 ? reg111[(1'h1):(1'h0)] : reg132);
  assign wire147 = reg117[(4'ha):(1'h1)];
  always
    @(posedge clk) begin
      reg148 <= ((~&$unsigned((!wire147))) >>> wire133);
      reg149 = ({$signed((reg129[(5'h13):(2'h3)] ? reg140 : (~reg139))),
              (reg130[(4'he):(3'h5)] ?
                  $signed(forvar110[(3'h7):(1'h0)]) : $unsigned((~&reg108)))} ?
          (-((7'h43) + ($unsigned(reg137) != (-reg130)))) : $signed(reg141[(1'h0):(1'h0)]));
    end
  assign wire150 = $unsigned(reg140[(1'h1):(1'h1)]);
  always
    @(posedge clk) begin
      reg151 <= (+((((reg149 ? wire145 : reg120) ?
              (8'hb7) : (reg111 ? reg138 : reg113)) ?
          $unsigned($signed(reg116)) : $unsigned(((8'hba) ~^ reg131))) <<< (((reg123 ?
              wire145 : reg144) >>> $unsigned((7'h43))) ?
          $signed(reg118[(4'h8):(1'h1)]) : (((8'ha4) != wire99) == reg106[(3'h4):(1'h0)]))));
      reg152 <= (~|reg130);
      reg153 = ({$signed(($signed(reg108) >= reg126[(2'h3):(1'h1)]))} ?
          reg108[(3'h7):(1'h1)] : $unsigned({reg123[(2'h3):(2'h3)]}));
      reg154 <= reg144;
    end
endmodule

module module39  (y, clk, wire44, wire43, wire42, wire41, wire40);
  output wire [(32'h196):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire44;
  input wire signed [(4'hb):(1'h0)] wire43;
  input wire signed [(5'h10):(1'h0)] wire42;
  input wire signed [(4'hf):(1'h0)] wire41;
  input wire [(4'hf):(1'h0)] wire40;
  wire signed [(4'hb):(1'h0)] wire77;
  wire signed [(4'he):(1'h0)] wire76;
  reg signed [(3'h4):(1'h0)] reg75 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg74 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg73 = (1'h0);
  reg [(5'h15):(1'h0)] reg72 = (1'h0);
  reg [(5'h12):(1'h0)] forvar71 = (1'h0);
  reg [(4'h9):(1'h0)] reg70 = (1'h0);
  reg [(4'he):(1'h0)] reg69 = (1'h0);
  reg [(5'h11):(1'h0)] reg68 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar67 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg66 = (1'h0);
  reg [(4'hd):(1'h0)] reg65 = (1'h0);
  reg [(4'hd):(1'h0)] reg64 = (1'h0);
  reg [(4'hb):(1'h0)] reg63 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg62 = (1'h0);
  reg [(5'h11):(1'h0)] reg61 = (1'h0);
  reg [(4'ha):(1'h0)] reg60 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg59 = (1'h0);
  reg [(3'h5):(1'h0)] reg58 = (1'h0);
  reg [(5'h12):(1'h0)] reg57 = (1'h0);
  reg [(4'h9):(1'h0)] reg56 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg55 = (1'h0);
  reg [(3'h4):(1'h0)] forvar54 = (1'h0);
  reg [(4'h9):(1'h0)] reg53 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar52 = (1'h0);
  reg [(4'hd):(1'h0)] reg51 = (1'h0);
  reg [(4'hc):(1'h0)] reg50 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg49 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg48 = (1'h0);
  reg [(4'ha):(1'h0)] reg47 = (1'h0);
  reg [(4'hc):(1'h0)] reg46 = (1'h0);
  wire [(5'h11):(1'h0)] wire45;
  assign y = {wire77,
                 wire76,
                 reg75,
                 reg74,
                 reg73,
                 reg72,
                 forvar71,
                 reg70,
                 reg69,
                 reg68,
                 forvar67,
                 reg66,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 reg55,
                 forvar54,
                 reg53,
                 forvar52,
                 reg51,
                 reg50,
                 reg49,
                 reg48,
                 reg47,
                 reg46,
                 wire45,
                 (1'h0)};
  assign wire45 = wire40;
  always
    @(posedge clk) begin
      reg46 <= wire40;
      reg47 <= wire40;
      reg48 <= $signed($signed((8'ha6)));
      reg49 = wire45;
    end
  always
    @(posedge clk) begin
      reg50 <= (-$unsigned(wire45));
      reg51 = ($signed((reg50 ~^ (wire40 ?
              ((8'hb3) < reg47) : (wire40 <= wire45)))) ?
          $signed({$unsigned((~|reg50)),
              (^~$signed(wire45))}) : $unsigned($signed(reg46[(3'h6):(3'h5)])));
      for (forvar52 = (1'h0); (forvar52 < (3'h4)); forvar52 = (forvar52 + (1'h1)))
        begin
          reg53 <= {((&(wire43 ?
                      ((7'h42) ? wire40 : wire44) : $signed(wire40))) ?
                  $unsigned(reg46[(3'h5):(2'h3)]) : wire41)};
          for (forvar54 = (1'h0); (forvar54 < (2'h2)); forvar54 = (forvar54 + (1'h1)))
            begin
              reg55 <= ((~|$unsigned(((reg49 ? forvar52 : reg48) ?
                      (8'hbe) : {wire45, reg50}))) ?
                  $unsigned((reg48[(4'ha):(2'h3)] + reg53)) : $signed(($unsigned(reg50) ?
                      (|forvar54[(3'h4):(2'h3)]) : (7'h43))));
              reg56 <= forvar52;
              reg57 <= wire42[(3'h4):(2'h2)];
              reg58 <= (|(wire40[(3'h6):(2'h2)] ?
                  $unsigned($unsigned($signed(wire44))) : ((|{forvar54}) > (reg57[(2'h2):(1'h1)] > $signed(reg48)))));
              reg59 <= (reg58[(1'h0):(1'h0)] ^~ ((+reg58[(3'h5):(2'h3)]) ?
                  reg47[(4'h8):(3'h5)] : (forvar54 ?
                      ($unsigned(wire43) == wire45) : (reg50[(4'h9):(2'h2)] ?
                          $unsigned(forvar52) : $signed(reg53)))));
            end
          reg60 <= (~|((($unsigned((8'hb6)) ?
                  reg55[(4'h9):(1'h0)] : $signed(forvar52)) != wire40) ?
              reg50[(3'h6):(1'h0)] : {{$signed(reg50), reg53[(3'h7):(3'h4)]},
                  (~|wire42[(3'h6):(2'h3)])}));
          reg61 = (!({{reg59[(2'h3):(2'h2)], ((8'hbe) >= reg53)}, wire44} ?
              (|reg53) : wire43[(4'h9):(4'h8)]));
          reg62 <= ((reg60 ?
              reg48[(5'h14):(2'h2)] : {$unsigned((^~reg56))}) == ({reg46,
                  reg53} ?
              $unsigned((|reg60[(3'h7):(1'h1)])) : (($signed((8'hb0)) ?
                  ((8'hb9) ?
                      reg59 : wire44) : reg46[(4'hb):(4'h8)]) ^ ((|wire42) ?
                  ((8'ha2) && (7'h40)) : (wire44 ? reg59 : (8'hb0))))));
        end
      reg63 <= $unsigned(wire42);
      reg64 <= $unsigned((($signed({wire44}) ?
          ($unsigned(reg59) << $signed((8'h9e))) : ((~^reg55) && $unsigned(wire43))) <<< wire42[(4'hc):(4'h8)]));
    end
  always
    @(posedge clk) begin
      reg65 <= ($signed(({(!wire44)} ^ reg53[(1'h0):(1'h0)])) && reg48[(4'h9):(2'h3)]);
      reg66 <= ((~|((~|(wire44 * (8'hb1))) ?
              $signed(reg50) : (-(wire42 && reg61)))) ?
          $unsigned(((&reg47[(1'h1):(1'h0)]) || ($unsigned(reg53) ?
              $signed(wire44) : reg60[(4'h9):(4'h9)]))) : (reg62[(4'h8):(3'h7)] & $unsigned(wire40)));
      for (forvar67 = (1'h0); (forvar67 < (2'h3)); forvar67 = (forvar67 + (1'h1)))
        begin
          reg68 <= $unsigned($unsigned(($signed(reg51[(4'hc):(2'h2)]) ^~ {{(8'hac),
                  wire45}})));
          reg69 <= ((reg58[(1'h1):(1'h0)] ?
              wire44[(4'h9):(3'h5)] : reg47) + reg57[(3'h4):(3'h4)]);
          reg70 = $unsigned((~^{(~^$unsigned((8'hbc))), {$unsigned(reg51)}}));
          for (forvar71 = (1'h0); (forvar71 < (1'h1)); forvar71 = (forvar71 + (1'h1)))
            begin
              reg72 <= ($unsigned(($unsigned(reg63) ?
                  $signed($unsigned(wire40)) : $unsigned($unsigned((8'h9e))))) != reg69);
              reg73 <= reg70;
            end
          reg74 <= reg51;
        end
      reg75 = $unsigned((reg73 ?
          ((reg66 | (^~reg66)) || ({forvar71} == reg58[(1'h1):(1'h1)])) : wire42));
    end
  assign wire76 = {$unsigned(wire42[(3'h7):(3'h6)])};
  assign wire77 = (reg50 < $signed($unsigned(reg73)));
endmodule

module module275
#( parameter param407 = {(~((^(|(8'hb7))) | ((&(8'ha2)) ? ((8'hb8) + (8'ha4)) : ((8'hba) ? (8'hb4) : (8'hb8))))), (~&(((~&(8'h9c)) ? ((8'h9e) ? (8'hac) : (8'ha2)) : ((8'had) ? (8'h9e) : (8'hb2))) < ({(8'haa)} ? ((8'h9e) >> (8'h9c)) : ((8'h9c) ? (8'hab) : (8'hb6)))))} )
(y, clk, wire279, wire278, wire277, wire276);
  output wire [(32'h200):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h9):(1'h0)] wire279;
  input wire signed [(2'h3):(1'h0)] wire278;
  input wire [(4'hb):(1'h0)] wire277;
  input wire signed [(3'h7):(1'h0)] wire276;
  reg [(5'h11):(1'h0)] reg406 = (1'h0);
  reg [(2'h2):(1'h0)] reg405 = (1'h0);
  reg [(4'h8):(1'h0)] reg404 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg403 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg402 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg401 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg400 = (1'h0);
  reg [(4'hc):(1'h0)] reg399 = (1'h0);
  reg [(5'h10):(1'h0)] reg398 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg397 = (1'h0);
  reg [(4'h9):(1'h0)] reg396 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar395 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar394 = (1'h0);
  reg [(3'h7):(1'h0)] reg393 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg392 = (1'h0);
  wire [(4'h9):(1'h0)] wire391;
  wire signed [(4'hb):(1'h0)] wire390;
  reg [(4'h8):(1'h0)] reg389 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg388 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg387 = (1'h0);
  reg [(3'h4):(1'h0)] reg386 = (1'h0);
  reg [(5'h14):(1'h0)] reg385 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire384;
  wire [(4'hc):(1'h0)] wire382;
  reg signed [(4'h8):(1'h0)] reg299 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg298 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg297 = (1'h0);
  reg [(4'ha):(1'h0)] reg296 = (1'h0);
  reg [(2'h3):(1'h0)] reg295 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar294 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire293;
  wire signed [(2'h2):(1'h0)] wire292;
  reg [(4'h8):(1'h0)] reg291 = (1'h0);
  reg [(4'hf):(1'h0)] reg290 = (1'h0);
  reg [(3'h5):(1'h0)] reg289 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg288 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg287 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar286 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg285 = (1'h0);
  reg [(4'hc):(1'h0)] reg284 = (1'h0);
  reg [(3'h6):(1'h0)] reg283 = (1'h0);
  reg [(2'h2):(1'h0)] reg282 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg281 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg280 = (1'h0);
  assign y = {reg406,
                 reg405,
                 reg404,
                 reg403,
                 reg402,
                 reg401,
                 reg400,
                 reg399,
                 reg398,
                 reg397,
                 reg396,
                 forvar395,
                 forvar394,
                 reg393,
                 reg392,
                 wire391,
                 wire390,
                 reg389,
                 reg388,
                 reg387,
                 reg386,
                 reg385,
                 wire384,
                 wire382,
                 reg299,
                 reg298,
                 reg297,
                 reg296,
                 reg295,
                 forvar294,
                 wire293,
                 wire292,
                 reg291,
                 reg290,
                 reg289,
                 reg288,
                 reg287,
                 forvar286,
                 reg285,
                 reg284,
                 reg283,
                 reg282,
                 reg281,
                 reg280,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg280 <= ($unsigned({wire279[(1'h0):(1'h0)]}) ?
          wire276 : $unsigned($unsigned($unsigned(wire278[(2'h3):(1'h1)]))));
      reg281 <= $signed($signed((($unsigned(wire278) ? (~|wire277) : wire278) ?
          {(wire279 | wire276)} : wire278)));
      reg282 <= (wire277 ? wire276 : (8'h9f));
    end
  always
    @(posedge clk) begin
      reg283 <= reg282[(1'h1):(1'h1)];
      reg284 <= ((+(wire276[(1'h1):(1'h0)] != $signed($signed((8'hab))))) ?
          ($signed((~^reg282[(1'h1):(1'h1)])) ^~ reg280[(3'h7):(3'h7)]) : wire277[(1'h1):(1'h0)]);
      reg285 <= (({$unsigned((reg283 && reg281)), $unsigned((+reg281))} ?
              (~|wire276[(3'h4):(1'h1)]) : wire278[(1'h0):(1'h0)]) ?
          $unsigned(wire279) : $unsigned(reg280[(4'hd):(4'h9)]));
    end
  always
    @(posedge clk) begin
      for (forvar286 = (1'h0); (forvar286 < (1'h0)); forvar286 = (forvar286 + (1'h1)))
        begin
          reg287 = $unsigned((~$signed((^~reg285[(4'hf):(4'h8)]))));
        end
      reg288 <= (-reg281);
      reg289 <= {((&(wire279 >= (forvar286 == reg280))) ?
              (|{forvar286[(4'he):(3'h7)]}) : forvar286)};
      reg290 <= (!wire276[(2'h3):(1'h0)]);
      reg291 <= ({reg290[(1'h1):(1'h1)]} ?
          ($unsigned(wire276) ^~ (reg284[(2'h3):(2'h2)] ?
              ($signed(wire278) ?
                  reg284[(3'h5):(2'h2)] : (wire277 ?
                      reg287 : wire279)) : reg280[(2'h3):(1'h1)])) : $unsigned(wire276[(2'h3):(2'h3)]));
    end
  assign wire292 = ($signed(({$signed(reg290),
                       forvar286[(4'ha):(3'h6)]} ~^ (8'hb3))) && wire279[(4'h9):(1'h0)]);
  assign wire293 = ({$signed({reg281, {reg291, forvar286}}),
                       wire278} < $signed((reg291[(2'h2):(1'h0)] * (-$signed(reg285)))));
  always
    @(posedge clk) begin
      for (forvar294 = (1'h0); (forvar294 < (1'h1)); forvar294 = (forvar294 + (1'h1)))
        begin
          reg295 <= reg289;
          reg296 <= $signed($unsigned(($signed(wire276) | $unsigned(wire293[(4'h9):(2'h2)]))));
        end
      reg297 <= wire293[(1'h0):(1'h0)];
      reg298 = $unsigned($unsigned((wire279 <= $unsigned(reg289[(2'h2):(1'h0)]))));
      reg299 <= wire292;
    end
  module300 modinst383 (wire382, clk, reg291, reg285, reg296, reg281);
  assign wire384 = ((~^((reg280 && (+(8'hb3))) ?
                       (((8'h9e) ^ (8'hbd)) ?
                           {(8'ha6)} : $signed((8'hab))) : (wire276[(3'h5):(3'h4)] >>> {forvar286}))) != {$unsigned((reg289[(3'h5):(2'h2)] ^~ {(8'hbb)})),
                       (8'hbd)});
  always
    @(posedge clk) begin
      reg385 <= ($signed($signed($signed((&reg280)))) - (($signed(reg284) ^~ reg289[(3'h5):(3'h4)]) != $unsigned(((~&reg298) != $signed(reg280)))));
      reg386 <= (+((+reg295) ?
          $unsigned($unsigned(reg290)) : reg298[(4'ha):(3'h6)]));
    end
  always
    @(posedge clk) begin
      reg387 <= ({wire293[(4'hd):(4'hc)]} == reg284);
      reg388 <= (&$signed(reg291[(1'h1):(1'h0)]));
      reg389 <= $unsigned(((((wire277 | wire277) ?
                  $unsigned(reg283) : (~|reg298)) ?
              (!reg386[(1'h0):(1'h0)]) : reg289) ?
          reg297[(4'hb):(1'h1)] : $signed($unsigned(reg282[(1'h0):(1'h0)]))));
    end
  assign wire390 = ((-$unsigned(reg289)) + ({(8'ha0)} ?
                       $unsigned(reg387) : {(reg297[(4'hd):(2'h3)] ?
                               reg285[(1'h1):(1'h0)] : (reg290 >> reg280)),
                           (reg288 ?
                               (reg385 ?
                                   wire382 : forvar286) : $unsigned(reg297))}));
  assign wire391 = wire279[(4'h9):(4'h8)];
  always
    @(posedge clk) begin
      reg392 <= wire382;
      reg393 <= ((~^(|((reg295 ? reg290 : reg283) ?
              $unsigned(reg385) : $signed((8'hb5))))) ?
          $signed(reg389[(3'h4):(1'h1)]) : wire391);
    end
  always
    @(posedge clk) begin
      for (forvar394 = (1'h0); (forvar394 < (3'h4)); forvar394 = (forvar394 + (1'h1)))
        begin
          for (forvar395 = (1'h0); (forvar395 < (1'h0)); forvar395 = (forvar395 + (1'h1)))
            begin
              reg396 = (!(~^(!{reg291, (reg389 | reg388)})));
              reg397 <= $unsigned(wire391[(4'h8):(3'h7)]);
              reg398 = ($unsigned(((+(wire390 ^ reg393)) ?
                  $signed($unsigned((7'h40))) : $signed((~reg288)))) > $unsigned(forvar294));
              reg399 = ({(^((reg299 * wire293) + {wire390, wire382})),
                      $signed($unsigned($signed(reg387)))} ?
                  forvar286 : reg282[(2'h2):(1'h0)]);
              reg400 <= reg397[(2'h2):(1'h0)];
            end
          reg401 <= $signed($signed(reg387[(3'h6):(2'h3)]));
          reg402 <= (^~$unsigned(reg284[(2'h2):(1'h0)]));
        end
      reg403 <= (~|forvar395[(3'h7):(3'h7)]);
      reg404 <= reg401[(4'hb):(3'h4)];
      reg405 <= ($unsigned(($signed((~&(8'hac))) ?
              wire391[(3'h5):(2'h3)] : $unsigned(reg388))) ?
          $unsigned($signed(reg289)) : $unsigned($unsigned((!reg399[(3'h6):(2'h2)]))));
      reg406 <= (forvar395 | (reg282[(2'h2):(2'h2)] ?
          wire279 : (reg402[(2'h2):(2'h2)] ?
              (reg299 - (wire391 == reg404)) : ({reg287,
                  wire278} || (^reg290)))));
    end
endmodule

module module231
#( parameter param258 = (((+(((8'h9e) == (8'haf)) ? ((8'hbe) ? (8'ha6) : (8'haa)) : (!(8'ha0)))) <<< (~^((~&(8'ha3)) ? {(8'h9e)} : ((8'hb9) >= (8'hbd))))) ? ((-(+(!(8'h9c)))) ? (+{(8'h9e)}) : {(((8'ha7) ^ (8'ha0)) ? (-(8'hb0)) : ((8'ha1) ^ (8'hbb))), (((8'hbd) || (7'h42)) && (-(8'h9e)))}) : ((({(8'hbe), (8'ha9)} ? ((8'h9e) ? (8'h9c) : (8'haf)) : ((8'hb0) ? (8'hb5) : (8'had))) ? (!(^~(8'hbd))) : (((8'ha5) ? (8'h9e) : (8'ha3)) ? (8'ha7) : ((8'hb6) ? (8'hbf) : (7'h40)))) ? ((8'hac) ^~ {{(8'hb0)}}) : {(~{(7'h41), (8'h9f)}), {((8'hb3) * (7'h44))}})) )
(y, clk, wire236, wire235, wire234, wire233, wire232);
  output wire [(32'hef):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'he):(1'h0)] wire236;
  input wire signed [(2'h3):(1'h0)] wire235;
  input wire signed [(4'hf):(1'h0)] wire234;
  input wire [(4'hf):(1'h0)] wire233;
  input wire [(3'h7):(1'h0)] wire232;
  reg signed [(3'h5):(1'h0)] reg257 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg256 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg255 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg254 = (1'h0);
  reg [(5'h10):(1'h0)] forvar253 = (1'h0);
  wire [(3'h6):(1'h0)] wire252;
  wire signed [(4'h8):(1'h0)] wire251;
  reg signed [(4'h9):(1'h0)] reg250 = (1'h0);
  reg [(5'h10):(1'h0)] reg249 = (1'h0);
  reg [(3'h7):(1'h0)] reg248 = (1'h0);
  reg [(5'h15):(1'h0)] reg247 = (1'h0);
  reg [(5'h11):(1'h0)] reg246 = (1'h0);
  reg [(3'h7):(1'h0)] reg245 = (1'h0);
  reg [(4'hf):(1'h0)] reg244 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg243 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg242 = (1'h0);
  reg [(5'h12):(1'h0)] reg241 = (1'h0);
  reg [(2'h3):(1'h0)] reg240 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar239 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar238 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg237 = (1'h0);
  assign y = {reg257,
                 reg256,
                 reg255,
                 reg254,
                 forvar253,
                 wire252,
                 wire251,
                 reg250,
                 reg249,
                 reg248,
                 reg247,
                 reg246,
                 reg245,
                 reg244,
                 reg243,
                 reg242,
                 reg241,
                 reg240,
                 forvar239,
                 forvar238,
                 reg237,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg237 <= $unsigned(($unsigned((~|(|wire236))) - (~|wire232[(2'h3):(2'h2)])));
      for (forvar238 = (1'h0); (forvar238 < (3'h4)); forvar238 = (forvar238 + (1'h1)))
        begin
          for (forvar239 = (1'h0); (forvar239 < (1'h1)); forvar239 = (forvar239 + (1'h1)))
            begin
              reg240 <= $unsigned({wire234[(3'h5):(3'h5)]});
              reg241 <= (((((+reg237) == (wire232 << reg237)) ?
                  (+wire236[(4'hc):(4'hc)]) : (|(wire234 + (8'haf)))) >> $signed($unsigned(((7'h43) <<< wire232)))) <<< wire233);
            end
          reg242 <= $unsigned($signed(reg237[(3'h5):(2'h3)]));
          if ((|reg240))
            begin
              reg243 = {wire232, wire233[(4'h8):(1'h0)]};
              reg244 <= (8'hbb);
              reg245 <= wire234;
              reg246 = $unsigned((~(((reg245 ?
                  wire233 : wire234) >> (reg244 ^ reg241)) << (!wire233[(4'hc):(4'hb)]))));
              reg247 <= (($unsigned(((!reg246) ?
                          ((8'hb6) || wire235) : $signed(wire232))) ?
                      ($signed((wire236 ? (8'hbe) : reg244)) ?
                          reg240[(1'h1):(1'h1)] : $signed((~|wire236))) : $unsigned($signed(forvar238[(3'h4):(3'h4)]))) ?
                  reg246[(4'h8):(3'h7)] : $signed(((^(|wire236)) << ((8'ha4) ?
                      (~^wire234) : $signed((8'hab))))));
            end
          else
            begin
              reg243 <= $unsigned((~$unsigned({forvar238, forvar239})));
              reg244 <= {$signed(wire236[(4'h8):(1'h1)]),
                  (-($signed((8'hb7)) != (~|{reg243, (8'hbb)})))};
              reg245 <= ((+$signed(((wire236 <= reg247) ?
                      $signed(wire232) : $unsigned(reg246)))) ?
                  (((wire234 == {reg240}) <= reg247) ?
                      ($unsigned(forvar239) >= (8'hbe)) : {reg246[(3'h7):(3'h4)]}) : (!($signed($unsigned(reg246)) ?
                      (8'ha5) : $signed((reg240 ? (8'ha9) : reg240)))));
            end
          reg248 <= $signed($unsigned(forvar239[(2'h2):(1'h1)]));
          reg249 <= reg243;
        end
      reg250 = ($unsigned($signed(wire233[(4'ha):(2'h2)])) == $unsigned(({{(8'hb5)},
              $unsigned(reg240)} ?
          reg244 : (^{wire235, reg247}))));
    end
  assign wire251 = ((^(-$unsigned($unsigned(reg240)))) != reg246);
  assign wire252 = $unsigned($unsigned($unsigned($signed($unsigned(reg243)))));
  always
    @(posedge clk) begin
      for (forvar253 = (1'h0); (forvar253 < (1'h1)); forvar253 = (forvar253 + (1'h1)))
        begin
          reg254 <= (forvar239[(2'h3):(2'h2)] ?
              $unsigned((((reg244 ^ wire252) != (^forvar239)) << wire234[(3'h5):(3'h4)])) : ((8'h9d) ?
                  (~^$unsigned($unsigned((8'ha9)))) : $signed({$signed(wire251)})));
          reg255 <= {(~|$unsigned(reg246))};
          reg256 <= $unsigned(wire252[(3'h5):(1'h1)]);
        end
      reg257 <= (wire235 ?
          wire252[(1'h1):(1'h1)] : (^~$signed(((8'hbf) >> (reg242 <= (8'hb5))))));
    end
endmodule

module module300
#( parameter param381 = (~{(!(((8'hbc) ? (7'h43) : (8'ha0)) + ((8'ha5) ^ (8'ha3)))), (8'ha5)}) )
(y, clk, wire304, wire303, wire302, wire301);
  output wire [(32'h16f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h6):(1'h0)] wire304;
  input wire signed [(4'h9):(1'h0)] wire303;
  input wire [(4'ha):(1'h0)] wire302;
  input wire signed [(4'hc):(1'h0)] wire301;
  reg [(4'ha):(1'h0)] reg380 = (1'h0);
  reg [(2'h3):(1'h0)] forvar379 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg378 = (1'h0);
  reg [(5'h12):(1'h0)] reg377 = (1'h0);
  wire [(5'h12):(1'h0)] wire376;
  wire signed [(3'h4):(1'h0)] wire374;
  wire signed [(3'h6):(1'h0)] wire328;
  reg [(5'h15):(1'h0)] reg327 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg326 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg325 = (1'h0);
  reg [(4'hb):(1'h0)] reg324 = (1'h0);
  reg [(5'h14):(1'h0)] forvar323 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg322 = (1'h0);
  reg [(3'h4):(1'h0)] reg321 = (1'h0);
  reg [(4'hb):(1'h0)] reg320 = (1'h0);
  reg [(3'h7):(1'h0)] reg319 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar318 = (1'h0);
  reg [(2'h2):(1'h0)] reg317 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire316;
  reg signed [(4'h9):(1'h0)] reg315 = (1'h0);
  reg [(3'h5):(1'h0)] reg314 = (1'h0);
  reg [(4'hd):(1'h0)] reg313 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg312 = (1'h0);
  reg [(4'h9):(1'h0)] reg311 = (1'h0);
  reg [(5'h11):(1'h0)] forvar310 = (1'h0);
  reg [(5'h12):(1'h0)] reg309 = (1'h0);
  reg [(2'h2):(1'h0)] reg308 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar307 = (1'h0);
  reg [(4'hc):(1'h0)] reg306 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire305;
  assign y = {reg380,
                 forvar379,
                 reg378,
                 reg377,
                 wire376,
                 wire374,
                 wire328,
                 reg327,
                 reg326,
                 reg325,
                 reg324,
                 forvar323,
                 reg322,
                 reg321,
                 reg320,
                 reg319,
                 forvar318,
                 reg317,
                 wire316,
                 reg315,
                 reg314,
                 reg313,
                 reg312,
                 reg311,
                 forvar310,
                 reg309,
                 reg308,
                 forvar307,
                 reg306,
                 wire305,
                 (1'h0)};
  assign wire305 = (^~wire301);
  always
    @(posedge clk) begin
      reg306 <= (^~wire301);
      for (forvar307 = (1'h0); (forvar307 < (2'h3)); forvar307 = (forvar307 + (1'h1)))
        begin
          reg308 = {((((wire302 ? wire302 : wire305) ?
                      (^wire302) : wire302[(1'h0):(1'h0)]) ?
                  (~&wire305) : (+(~&forvar307))) >> reg306[(4'hc):(4'h9)])};
          reg309 <= $signed(forvar307);
          for (forvar310 = (1'h0); (forvar310 < (1'h1)); forvar310 = (forvar310 + (1'h1)))
            begin
              reg311 = reg308[(1'h1):(1'h1)];
              reg312 = $signed($signed((~|$signed(wire302))));
              reg313 <= ({{reg311, wire304}, $signed(reg306)} ^ (8'haf));
              reg314 = reg309[(2'h3):(2'h2)];
            end
          reg315 <= $signed((((wire305[(1'h1):(1'h1)] != forvar310[(3'h4):(1'h0)]) ?
                  $unsigned((8'hbe)) : $signed($unsigned(reg312))) ?
              (|(+(reg308 ? reg313 : reg306))) : wire303[(3'h5):(1'h0)]));
        end
    end
  assign wire316 = $signed(((((wire305 && (8'hb7)) + (8'hbb)) != forvar310) ^ $signed(forvar310[(4'hb):(3'h5)])));
  always
    @(posedge clk) begin
      reg317 <= wire302;
      for (forvar318 = (1'h0); (forvar318 < (2'h2)); forvar318 = (forvar318 + (1'h1)))
        begin
          reg319 <= (wire304[(1'h1):(1'h0)] <<< ($unsigned(reg315) ?
              wire316[(1'h0):(1'h0)] : ($signed($unsigned(forvar307)) << $unsigned($signed(reg309)))));
          reg320 = forvar318[(5'h12):(5'h12)];
          reg321 <= ($unsigned((($unsigned(wire303) ?
              $unsigned(reg320) : (forvar310 || wire305)) < $signed((reg306 ?
              (8'hb2) : reg314)))) > (8'h9c));
        end
    end
  always
    @(posedge clk) begin
      reg322 <= (reg313 || $signed(wire316));
      for (forvar323 = (1'h0); (forvar323 < (2'h3)); forvar323 = (forvar323 + (1'h1)))
        begin
          reg324 <= ($signed((+wire305[(3'h4):(3'h4)])) + wire316);
          reg325 = wire301;
          reg326 <= (8'hb6);
        end
      reg327 <= (wire316 ?
          reg308 : ({reg326} == {{(reg313 ? reg320 : (7'h42)),
                  $signed(reg320)}}));
    end
  assign wire328 = ($unsigned(reg306) != $unsigned(reg324[(4'h8):(1'h0)]));
  module329 modinst375 (wire374, clk, reg326, reg327, reg320, reg313);
  assign wire376 = {{reg311}, {{$signed(reg324)}}};
  always
    @(posedge clk) begin
      reg377 <= reg325;
      reg378 <= reg377;
      for (forvar379 = (1'h0); (forvar379 < (2'h3)); forvar379 = (forvar379 + (1'h1)))
        begin
          reg380 <= (&($unsigned((8'hac)) | (($signed(wire304) ?
              $unsigned(reg321) : wire305[(5'h10):(3'h4)]) <<< $signed((wire304 >> wire301)))));
        end
    end
endmodule

module module329
#( parameter param372 = (~&(|((+{(7'h41), (7'h42)}) ? (((8'ha6) != (8'h9c)) ? ((8'hb6) ? (8'ha2) : (8'hb2)) : ((8'hbd) ^ (8'h9d))) : (~^((8'hba) > (8'hac))))))
, parameter param373 = (param372 & (~|(((param372 > param372) == {param372, param372}) ? (!{(8'hb7), param372}) : ((8'hb2) ^ (param372 ? param372 : param372))))) )
(y, clk, wire333, wire332, wire331, wire330);
  output wire [(32'h205):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire333;
  input wire signed [(4'hd):(1'h0)] wire332;
  input wire signed [(3'h5):(1'h0)] wire331;
  input wire [(4'hd):(1'h0)] wire330;
  reg signed [(5'h11):(1'h0)] reg371 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg370 = (1'h0);
  reg [(2'h3):(1'h0)] reg369 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire368;
  wire signed [(4'hc):(1'h0)] wire367;
  reg [(5'h12):(1'h0)] reg366 = (1'h0);
  reg [(5'h15):(1'h0)] reg365 = (1'h0);
  reg [(4'hb):(1'h0)] reg364 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg363 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar362 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg361 = (1'h0);
  reg [(2'h3):(1'h0)] reg360 = (1'h0);
  reg [(2'h3):(1'h0)] forvar359 = (1'h0);
  reg [(5'h14):(1'h0)] reg358 = (1'h0);
  reg [(4'he):(1'h0)] reg357 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar356 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg355 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg354 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg353 = (1'h0);
  reg [(5'h10):(1'h0)] reg352 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg351 = (1'h0);
  reg [(4'ha):(1'h0)] forvar350 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg349 = (1'h0);
  reg [(5'h11):(1'h0)] reg348 = (1'h0);
  wire [(5'h15):(1'h0)] wire347;
  wire [(5'h13):(1'h0)] wire346;
  wire [(4'hd):(1'h0)] wire345;
  reg signed [(5'h10):(1'h0)] reg344 = (1'h0);
  wire [(5'h15):(1'h0)] wire343;
  reg signed [(5'h14):(1'h0)] reg342 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg341 = (1'h0);
  reg [(5'h13):(1'h0)] reg340 = (1'h0);
  reg [(3'h4):(1'h0)] reg339 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar338 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg337 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg336 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg335 = (1'h0);
  reg [(4'hf):(1'h0)] reg334 = (1'h0);
  assign y = {reg371,
                 reg370,
                 reg369,
                 wire368,
                 wire367,
                 reg366,
                 reg365,
                 reg364,
                 reg363,
                 forvar362,
                 reg361,
                 reg360,
                 forvar359,
                 reg358,
                 reg357,
                 forvar356,
                 reg355,
                 reg354,
                 reg353,
                 reg352,
                 reg351,
                 forvar350,
                 reg349,
                 reg348,
                 wire347,
                 wire346,
                 wire345,
                 reg344,
                 wire343,
                 reg342,
                 reg341,
                 reg340,
                 reg339,
                 forvar338,
                 reg337,
                 reg336,
                 reg335,
                 reg334,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg334 = (wire332 ?
          $unsigned(wire333) : (((wire331[(1'h1):(1'h0)] ?
              (8'hb6) : (8'hb7)) * ((wire332 ? wire330 : wire331) ?
              (~&wire331) : (wire330 ? wire332 : wire333))) == (8'hb5)));
      reg335 <= wire333[(2'h2):(1'h0)];
      reg336 = (8'hb2);
    end
  always
    @(posedge clk) begin
      reg337 = ($signed((^~(wire332 + $unsigned(reg334)))) ^~ $signed($signed(reg336)));
      for (forvar338 = (1'h0); (forvar338 < (3'h4)); forvar338 = (forvar338 + (1'h1)))
        begin
          reg339 <= $unsigned({$unsigned(reg336[(3'h4):(1'h1)])});
        end
      reg340 = (({wire333} ?
              wire332[(4'h9):(3'h5)] : $unsigned($unsigned((!wire332)))) ?
          (reg339[(2'h2):(1'h0)] <= ($signed(((8'hb4) ? reg337 : wire330)) ?
              (reg334 ^~ reg339[(1'h0):(1'h0)]) : (reg337[(4'h9):(2'h2)] ?
                  (~(8'h9f)) : ((8'ha6) >> reg334)))) : $unsigned(((~&$signed(reg336)) ?
              reg335 : $signed(wire333[(4'hf):(4'h9)]))));
      reg341 <= reg340;
      reg342 <= (~&($signed(reg335[(3'h5):(3'h5)]) ?
          $unsigned(((~^reg337) <<< (8'haa))) : $signed(reg334[(3'h5):(2'h2)])));
    end
  assign wire343 = (($signed(reg341[(3'h4):(2'h2)]) != (((wire332 <= wire332) && ((8'hb2) | wire333)) == reg334[(3'h6):(3'h6)])) != (^(8'ha6)));
  always
    @(posedge clk) begin
      reg344 = ({reg341, (&reg340)} == $signed((wire343 >> reg341)));
    end
  assign wire345 = (((reg341[(5'h10):(4'hf)] ?
                       $unsigned(reg337[(4'h9):(4'h8)]) : (+reg341[(4'ha):(1'h0)])) >>> $unsigned({(~reg341)})) <<< {$unsigned({reg335[(5'h12):(1'h0)],
                           reg340})});
  assign wire346 = $signed((|(~|{$signed(reg339), $unsigned((8'ha8))})));
  assign wire347 = $signed(wire331[(3'h5):(3'h5)]);
  always
    @(posedge clk) begin
      reg348 <= reg340;
      reg349 <= (~&(wire347 ~^ reg335));
      for (forvar350 = (1'h0); (forvar350 < (2'h3)); forvar350 = (forvar350 + (1'h1)))
        begin
          reg351 <= {(|reg348), wire346[(4'hb):(3'h4)]};
          reg352 <= wire346;
        end
      reg353 = wire347;
    end
  always
    @(posedge clk) begin
      reg354 <= ($signed((8'h9f)) ?
          ($signed({$unsigned(wire330)}) || wire343) : reg348);
      reg355 <= (~&((reg352 ?
          $signed((reg335 || wire331)) : $unsigned((reg349 ?
              wire330 : reg349))) == reg352[(4'hd):(4'hd)]));
      for (forvar356 = (1'h0); (forvar356 < (1'h1)); forvar356 = (forvar356 + (1'h1)))
        begin
          reg357 <= $signed((8'hac));
          reg358 <= {wire347[(1'h1):(1'h0)]};
        end
      for (forvar359 = (1'h0); (forvar359 < (2'h2)); forvar359 = (forvar359 + (1'h1)))
        begin
          reg360 <= reg352;
          reg361 <= $unsigned(((^~((reg344 & reg334) >>> (reg337 ?
              (8'hae) : wire331))) ^ wire332));
          for (forvar362 = (1'h0); (forvar362 < (3'h4)); forvar362 = (forvar362 + (1'h1)))
            begin
              reg363 <= {(^~reg334)};
              reg364 <= {($signed(reg349[(3'h5):(3'h4)]) | reg349[(3'h5):(2'h3)])};
              reg365 <= ({(~($unsigned(reg340) && (wire343 + wire343))),
                  ($unsigned((reg337 ? (8'hbb) : forvar356)) ?
                      (wire332 ?
                          $signed(reg364) : ((8'hb6) <= reg339)) : {$signed(reg335)})} >= (8'hb8));
            end
        end
      reg366 <= $unsigned(forvar359[(2'h3):(2'h2)]);
    end
  assign wire367 = (-reg349);
  assign wire368 = $signed((-forvar362));
  always
    @(posedge clk) begin
      reg369 <= $signed(reg341[(3'h5):(3'h5)]);
    end
  always
    @(posedge clk) begin
      reg370 <= reg361;
      reg371 <= (~^(|({$signed(reg364)} ?
          wire347[(4'he):(3'h7)] : reg342[(4'ha):(3'h6)])));
    end
endmodule