(* use_dsp48="no" *) (* use_dsp="no" *) module top
#( parameter param338 = {(8'hb8)}
, parameter param339 = ((~&(~&((param338 + param338) ? (param338 ? param338 : (8'h9f)) : param338))) ? (8'hba) : (({param338} <<< (+(~^param338))) <= (+{(param338 < param338), (^~param338)}))) )
(y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h37f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire0;
  input wire [(2'h2):(1'h0)] wire1;
  input wire signed [(5'h14):(1'h0)] wire2;
  input wire [(5'h10):(1'h0)] wire3;
  input wire [(4'hf):(1'h0)] wire4;
  reg [(5'h12):(1'h0)] reg337 = (1'h0);
  reg [(4'hd):(1'h0)] reg336 = (1'h0);
  reg signed [(4'he):(1'h0)] reg335 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg334 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg333 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg332 = (1'h0);
  reg [(3'h4):(1'h0)] reg331 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg330 = (1'h0);
  reg [(3'h4):(1'h0)] reg329 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg328 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg327 = (1'h0);
  wire [(4'ha):(1'h0)] wire326;
  wire [(3'h7):(1'h0)] wire324;
  wire signed [(4'h9):(1'h0)] wire197;
  wire [(4'hf):(1'h0)] wire5;
  wire [(4'h9):(1'h0)] wire6;
  reg signed [(3'h5):(1'h0)] reg7 = (1'h0);
  reg [(4'hf):(1'h0)] reg8 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg9 = (1'h0);
  reg [(4'he):(1'h0)] reg10 = (1'h0);
  reg [(4'hf):(1'h0)] reg11 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg12 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg13 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg14 = (1'h0);
  reg [(4'hd):(1'h0)] reg15 = (1'h0);
  reg [(3'h4):(1'h0)] reg16 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg17 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg18 = (1'h0);
  reg [(2'h2):(1'h0)] reg19 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg20 = (1'h0);
  reg [(4'h8):(1'h0)] reg21 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg22 = (1'h0);
  reg [(5'h11):(1'h0)] reg23 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg24 = (1'h0);
  reg [(2'h3):(1'h0)] reg25 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg26 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg27 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg28 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg29 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire30;
  wire signed [(4'h8):(1'h0)] wire31;
  wire signed [(3'h5):(1'h0)] wire32;
  wire [(5'h14):(1'h0)] wire33;
  wire [(4'ha):(1'h0)] wire34;
  wire signed [(5'h13):(1'h0)] wire35;
  reg [(4'hc):(1'h0)] reg36 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg37 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg38 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg39 = (1'h0);
  reg [(4'hf):(1'h0)] reg40 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg41 = (1'h0);
  reg [(2'h3):(1'h0)] reg42 = (1'h0);
  reg [(3'h4):(1'h0)] reg43 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg44 = (1'h0);
  reg [(5'h11):(1'h0)] reg45 = (1'h0);
  reg [(4'he):(1'h0)] reg46 = (1'h0);
  reg [(4'h9):(1'h0)] reg47 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg48 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg49 = (1'h0);
  reg [(3'h4):(1'h0)] reg50 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg51 = (1'h0);
  reg [(5'h10):(1'h0)] reg52 = (1'h0);
  reg [(3'h7):(1'h0)] reg53 = (1'h0);
  reg [(5'h14):(1'h0)] reg54 = (1'h0);
  reg [(5'h12):(1'h0)] reg55 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg56 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg57 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg58 = (1'h0);
  reg [(3'h6):(1'h0)] reg59 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg60 = (1'h0);
  reg [(4'h9):(1'h0)] reg61 = (1'h0);
  wire [(5'h12):(1'h0)] wire62;
  wire [(4'h9):(1'h0)] wire63;
  wire [(4'hb):(1'h0)] wire64;
  wire [(5'h11):(1'h0)] wire65;
  wire [(5'h12):(1'h0)] wire195;
  assign y = {reg337,
                 reg336,
                 reg335,
                 reg334,
                 reg333,
                 reg332,
                 reg331,
                 reg330,
                 reg329,
                 reg328,
                 reg327,
                 wire326,
                 wire324,
                 wire197,
                 wire5,
                 wire6,
                 reg7,
                 reg8,
                 reg9,
                 reg10,
                 reg11,
                 reg12,
                 reg13,
                 reg14,
                 reg15,
                 reg16,
                 reg17,
                 reg18,
                 reg19,
                 reg20,
                 reg21,
                 reg22,
                 reg23,
                 reg24,
                 reg25,
                 reg26,
                 reg27,
                 reg28,
                 reg29,
                 wire30,
                 wire31,
                 wire32,
                 wire33,
                 wire34,
                 wire35,
                 reg36,
                 reg37,
                 reg38,
                 reg39,
                 reg40,
                 reg41,
                 reg42,
                 reg43,
                 reg44,
                 reg45,
                 reg46,
                 reg47,
                 reg48,
                 reg49,
                 reg50,
                 reg51,
                 reg52,
                 reg53,
                 reg54,
                 reg55,
                 reg56,
                 reg57,
                 reg58,
                 reg59,
                 reg60,
                 reg61,
                 wire62,
                 wire63,
                 wire64,
                 wire65,
                 wire195,
                 (1'h0)};
  assign wire5 = $signed($signed((^{$signed(wire1), (wire2 - wire0)})));
  assign wire6 = wire5[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      if ($unsigned($unsigned($signed(wire6[(1'h1):(1'h1)]))))
        begin
          reg7 <= (^~(~$unsigned($signed(wire6[(3'h5):(1'h1)]))));
          reg8 <= $unsigned({wire4});
          if ((wire6 ~^ {wire3}))
            begin
              reg9 <= $unsigned($signed({wire2}));
              reg10 <= ($signed((($unsigned((8'hb9)) ?
                          wire4[(4'h8):(3'h5)] : $signed(wire1)) ?
                      wire3[(1'h1):(1'h0)] : (wire6 ^ $unsigned(reg9)))) ?
                  reg7[(1'h1):(1'h0)] : $signed((+(&wire5[(2'h2):(1'h1)]))));
              reg11 <= wire2;
              reg12 <= $signed($signed((~&$signed($unsigned(reg9)))));
            end
          else
            begin
              reg9 <= wire5[(3'h5):(1'h0)];
              reg10 <= $signed(reg10);
            end
          if (wire4[(4'h9):(2'h3)])
            begin
              reg13 <= reg7[(2'h3):(2'h3)];
              reg14 <= $signed((wire2[(2'h3):(1'h0)] > reg11[(4'h8):(2'h3)]));
              reg15 <= $signed(wire0);
              reg16 <= $unsigned({($unsigned($unsigned(reg7)) ?
                      $unsigned((reg10 ?
                          reg11 : wire0)) : ($unsigned(wire6) | wire4[(3'h7):(1'h0)])),
                  reg10});
              reg17 <= reg12[(4'hb):(4'hb)];
            end
          else
            begin
              reg13 <= wire1[(2'h2):(2'h2)];
              reg14 <= wire0;
              reg15 <= wire3;
              reg16 <= reg15[(2'h3):(1'h0)];
            end
        end
      else
        begin
          if ({((~|{$unsigned(wire3),
                  {wire0, (8'hbf)}}) >> ((~|$signed(reg11)) ?
                  (wire5[(4'ha):(3'h6)] - $unsigned(wire5)) : wire3))})
            begin
              reg7 <= (((wire4 >>> {$unsigned((8'haf)),
                      wire3[(4'h9):(4'h9)]}) ^ (((^reg15) ?
                      $signed((8'hb1)) : reg10[(4'h8):(3'h5)]) ^ wire0[(1'h0):(1'h0)])) ?
                  wire2[(5'h10):(5'h10)] : wire3);
              reg8 <= reg12[(4'hc):(4'h8)];
            end
          else
            begin
              reg7 <= $unsigned(reg15);
              reg8 <= (wire2[(3'h4):(2'h3)] > (~((8'hae) ?
                  ({reg9} ?
                      $signed(reg10) : reg7) : $signed($unsigned(reg12)))));
              reg9 <= (reg9[(3'h7):(3'h7)] ?
                  wire2 : (reg15 * reg15[(2'h2):(2'h2)]));
              reg10 <= (8'h9e);
              reg11 <= reg9[(4'hd):(4'h9)];
            end
          reg12 <= (!{({{reg9}, $unsigned(wire0)} ?
                  wire0[(3'h5):(1'h1)] : reg15),
              {((wire2 ? (8'ha6) : (8'hba)) ^ reg11), ((!reg16) && (^wire4))}});
        end
      reg18 <= wire1;
      if ((8'h9d))
        begin
          if (($signed({((^reg12) ? wire5 : {reg18, reg8})}) ?
              (~^($signed(wire6[(1'h0):(1'h0)]) * {$unsigned(reg13)})) : {(reg17[(3'h5):(3'h5)] | {reg11[(3'h6):(2'h3)],
                      {wire1, wire3}}),
                  (^($signed(reg16) ? wire6 : {wire3, reg13}))}))
            begin
              reg19 <= $signed(({$signed(wire6[(1'h0):(1'h0)])} ^ $unsigned(((8'hb5) && (reg13 && reg8)))));
              reg20 <= $signed(reg19);
              reg21 <= $signed({(wire5[(4'h9):(2'h2)] ?
                      $unsigned(((8'ha8) & wire0)) : (|$unsigned(reg17)))});
              reg22 <= wire2;
              reg23 <= ($unsigned(reg18[(3'h5):(2'h2)]) >> $signed($unsigned((|$signed((8'ha2))))));
            end
          else
            begin
              reg19 <= reg21;
              reg20 <= $unsigned($signed(($unsigned(((8'hb0) ~^ reg21)) ?
                  $unsigned(((8'ha4) ? reg23 : wire1)) : $signed((8'ha9)))));
              reg21 <= {{reg16[(2'h2):(2'h2)], $unsigned(reg17[(3'h4):(2'h2)])},
                  ($unsigned(reg10) ?
                      (reg7[(2'h2):(1'h1)] & (^$unsigned(reg18))) : $signed(wire1))};
            end
          reg24 <= $unsigned((7'h43));
          reg25 <= $signed(reg21[(1'h0):(1'h0)]);
          if ($signed((((~|(reg13 ? reg18 : wire5)) == (8'ha7)) ?
              {{{wire6, reg11}}} : (&(reg15[(3'h4):(3'h4)] ?
                  wire1 : reg9[(5'h11):(4'hd)])))))
            begin
              reg26 <= reg24;
            end
          else
            begin
              reg26 <= $unsigned(reg14);
              reg27 <= ({reg9[(3'h6):(2'h3)],
                  (wire6 | $signed(reg7[(1'h0):(1'h0)]))} >> ($signed($signed(reg23)) >>> reg22[(1'h1):(1'h1)]));
            end
        end
      else
        begin
          reg19 <= {((8'hbb) ?
                  (8'hb2) : {((~&reg17) ?
                          ((8'hbf) | reg11) : $unsigned((7'h41)))}),
              {($signed(((7'h43) ? (7'h43) : reg17)) ?
                      reg24 : ((|wire3) ? $signed((8'hbf)) : (reg17 && reg8))),
                  (~{(!(8'haa)), $signed(wire2)})}};
          reg20 <= $unsigned({reg8[(4'h8):(3'h7)],
              $signed({(reg20 ? wire5 : (8'ha2))})});
          reg21 <= (((((reg7 ? (8'hb6) : reg26) ?
                      reg17[(1'h0):(1'h0)] : {reg27,
                          wire0}) + $unsigned(wire5[(4'hf):(3'h5)])) ?
                  (7'h43) : reg13) ?
              ($unsigned({{reg16}, $signed(reg25)}) ?
                  $signed(reg20[(2'h2):(1'h0)]) : reg22[(2'h2):(1'h0)]) : (&($signed((wire0 > reg15)) ?
                  reg16[(3'h4):(1'h0)] : reg7)));
          reg22 <= wire0;
        end
      reg28 <= {$signed((($signed(reg14) ?
              (^~reg18) : (reg13 ~^ (8'hae))) >>> (reg22 <= (~|reg25)))),
          reg15[(2'h3):(2'h3)]};
      reg29 <= $signed(((!reg16) != $signed((wire0 ^ (wire3 ?
          (8'h9f) : wire5)))));
    end
  assign wire30 = reg26;
  assign wire31 = (($signed($signed($signed(reg8))) ?
                      {wire4[(4'hd):(3'h4)],
                          (reg21 ?
                              reg8 : $unsigned((8'hb5)))} : $signed(((8'hbf) || $unsigned(reg22)))) >= ((((reg13 == reg16) ?
                              (reg9 ? reg7 : reg24) : reg8[(2'h3):(2'h3)]) ?
                          (~^$signed(reg27)) : $signed($unsigned(reg18))) ?
                      $signed(wire6) : (^reg18)));
  assign wire32 = reg10;
  assign wire33 = ($signed(((8'hab) >>> reg20[(1'h0):(1'h0)])) ^ ({(-reg16)} && (~|((~wire3) && (^~reg9)))));
  assign wire34 = $signed($unsigned(reg11));
  assign wire35 = reg15[(3'h7):(2'h2)];
  always
    @(posedge clk) begin
      reg36 <= (~wire1[(1'h0):(1'h0)]);
      if (((!$signed(reg36[(2'h3):(2'h3)])) > (|reg16[(2'h3):(1'h0)])))
        begin
          reg37 <= reg13;
        end
      else
        begin
          reg37 <= reg10[(2'h3):(1'h1)];
          reg38 <= (^((($unsigned(reg23) <<< (wire2 ? wire3 : wire6)) ?
              $unsigned((reg29 > reg22)) : reg19[(1'h0):(1'h0)]) - ((reg29 & (!(8'ha5))) ?
              reg10[(4'hb):(1'h1)] : $signed(reg13[(1'h0):(1'h0)]))));
          reg39 <= ((8'ha3) ? $signed($signed({$unsigned(reg27)})) : reg19);
        end
    end
  always
    @(posedge clk) begin
      if (((reg10[(2'h2):(2'h2)] ? reg17 : reg9) - reg21[(2'h2):(2'h2)]))
        begin
          reg40 <= {$signed($unsigned(($signed((8'hba)) ?
                  (reg26 ? wire2 : (7'h43)) : (wire2 ? wire35 : wire0)))),
              $signed((reg17[(2'h3):(2'h3)] >= wire2[(5'h14):(4'hc)]))};
          reg41 <= (|reg11[(3'h7):(3'h4)]);
          reg42 <= ((~$signed(((reg11 <<< reg13) ~^ reg23[(3'h5):(2'h3)]))) ?
              wire2[(4'hf):(3'h6)] : $unsigned($signed((~&(!wire33)))));
        end
      else
        begin
          reg40 <= $unsigned($unsigned((reg9[(4'he):(4'ha)] ?
              ($signed(reg19) ?
                  (reg10 >= reg27) : (reg29 ?
                      reg19 : (8'hb6))) : reg13[(1'h1):(1'h0)])));
          reg41 <= (reg23[(4'hd):(4'hc)] * $unsigned((wire3[(1'h0):(1'h0)] == wire35[(4'he):(3'h6)])));
        end
    end
  always
    @(posedge clk) begin
      if (reg24)
        begin
          if ($unsigned(reg16[(2'h2):(1'h0)]))
            begin
              reg43 <= ($unsigned((($unsigned(wire35) ?
                      $signed(reg14) : ((8'ha9) ?
                          wire2 : wire34)) - ({reg38} == (|reg27)))) ?
                  wire2 : wire35[(4'h9):(3'h7)]);
              reg44 <= (({{(reg26 ? reg36 : wire1)},
                      wire2[(3'h7):(3'h7)]} || $signed(($unsigned((8'hb1)) ?
                      $unsigned(wire3) : ((8'hb4) ? wire0 : reg19)))) ?
                  ($signed(wire33) >>> (~(reg43 << (&wire4)))) : reg43[(2'h3):(2'h3)]);
            end
          else
            begin
              reg43 <= wire30[(5'h12):(4'hf)];
            end
          if ((8'ha1))
            begin
              reg45 <= (reg9[(3'h7):(1'h0)] ?
                  {{reg39}, wire0} : reg39[(3'h7):(3'h5)]);
              reg46 <= (~^(8'hbd));
              reg47 <= {reg24[(4'hb):(3'h6)],
                  $unsigned((-$signed((wire0 ? wire1 : reg18))))};
            end
          else
            begin
              reg45 <= reg25[(1'h0):(1'h0)];
              reg46 <= (!(&$signed({$signed(reg27)})));
            end
          reg48 <= {reg38[(3'h6):(1'h0)], (8'hbe)};
          reg49 <= $signed(reg47);
        end
      else
        begin
          if ($unsigned((|(^~$unsigned($unsigned(reg23))))))
            begin
              reg43 <= reg21;
            end
          else
            begin
              reg43 <= ($signed(reg24) && $unsigned((({reg14} + (reg28 >= (8'ha9))) ^ $unsigned((~|(8'ha0))))));
              reg44 <= ({reg45[(4'hc):(1'h0)]} && $signed((($unsigned(reg14) ?
                      (~&(8'ha9)) : $signed(reg46)) ?
                  ((reg7 ~^ reg37) ~^ $signed(reg27)) : $signed($unsigned(reg25)))));
              reg45 <= reg37;
              reg46 <= (($signed($signed(((8'hb7) + wire32))) + $signed(reg9)) ?
                  reg48[(2'h2):(1'h1)] : (8'hac));
            end
          if ((~|(^~((8'ha3) >= $unsigned(reg20)))))
            begin
              reg47 <= reg28[(4'he):(4'hd)];
              reg48 <= ($signed(wire5) ?
                  ($signed(($unsigned(reg13) && {wire4,
                      reg44})) <<< $unsigned(reg46)) : ((((reg17 ?
                          wire35 : reg45) ?
                      (reg43 ?
                          (8'hba) : reg8) : reg47[(1'h0):(1'h0)]) >> $signed(reg9)) + reg28));
              reg49 <= {$unsigned((~^((!reg44) << (|reg38)))), (-(8'hae))};
            end
          else
            begin
              reg47 <= (^((~|(reg7[(2'h2):(1'h0)] ?
                  (8'hbc) : $unsigned((8'hb0)))) ^~ reg23));
              reg48 <= ((($unsigned(wire1) ?
                          reg40[(4'he):(4'hc)] : (wire3 >> reg43[(1'h1):(1'h0)])) ?
                      (((reg29 || reg27) ?
                          (reg49 * (8'hbc)) : reg26[(2'h2):(1'h0)]) * $unsigned(reg40[(3'h5):(2'h2)])) : ((((8'h9c) ?
                          reg10 : reg36) | wire31[(1'h0):(1'h0)]) != ((~^reg16) ?
                          (reg36 * reg16) : (|reg49)))) ?
                  wire5[(2'h3):(1'h1)] : (+reg21[(4'h8):(2'h3)]));
              reg49 <= {$signed($signed((8'h9e))),
                  (({(reg9 >>> reg29)} * (&(|reg36))) == reg24[(2'h3):(1'h1)])};
              reg50 <= (~(wire32[(1'h0):(1'h0)] < $unsigned($signed(reg36[(4'ha):(4'h9)]))));
              reg51 <= (wire33 <<< wire4[(2'h3):(1'h1)]);
            end
          reg52 <= reg9[(5'h10):(4'hb)];
          reg53 <= reg48;
        end
      reg54 <= $unsigned((!$signed(((^~wire5) ?
          $unsigned(reg49) : reg52[(4'hb):(3'h6)]))));
      reg55 <= (reg49[(4'hc):(1'h1)] ?
          reg27 : (wire3 ? (&(((8'ha1) | reg15) ? {wire3} : wire2)) : reg14));
      if (reg9)
        begin
          reg56 <= $signed(reg11);
          reg57 <= reg42[(2'h2):(1'h1)];
          reg58 <= (($signed({(^(8'hba)), {reg43, reg56}}) ?
              (-$signed($signed(reg11))) : (+(|$signed(wire34)))) | reg43[(2'h2):(1'h0)]);
          reg59 <= ((reg55[(4'hc):(1'h1)] && $signed(reg49)) >> reg14);
          reg60 <= $signed((!wire30));
        end
      else
        begin
          reg56 <= reg59[(1'h0):(1'h0)];
          reg57 <= wire0[(4'hc):(3'h4)];
          reg58 <= {reg23};
          reg59 <= reg11;
        end
      reg61 <= $signed((reg42 <= $unsigned(($unsigned((8'had)) == reg43))));
    end
  assign wire62 = (|($signed($signed((reg7 ? reg10 : (8'haa)))) ?
                      (reg46[(2'h3):(2'h2)] ?
                          (reg60[(1'h0):(1'h0)] * {(7'h40)}) : {(wire3 > reg13),
                              wire33}) : ($signed((reg38 | reg52)) != $unsigned(reg37[(2'h2):(1'h1)]))));
  assign wire63 = (^(&reg7));
  assign wire64 = (reg37 > reg60);
  assign wire65 = $unsigned((-reg17[(3'h4):(2'h2)]));
  module66 modinst196 (.wire68(reg15), .wire70(reg40), .wire71(reg55), .wire67(reg27), .y(wire195), .clk(clk), .wire69(wire64));
  assign wire197 = ($signed((((reg57 >>> reg44) ?
                           $unsigned(reg59) : reg41) + $signed(reg37))) ?
                       $unsigned(($signed((wire0 <= reg9)) ^~ $signed(((7'h42) ?
                           reg13 : reg49)))) : ($unsigned(reg47[(1'h0):(1'h0)]) + reg27));
  module198 modinst325 (wire324, clk, wire65, reg45, reg56, wire2);
  assign wire326 = (8'ha2);
  always
    @(posedge clk) begin
      if ($unsigned((8'had)))
        begin
          reg327 <= (^{wire1, $unsigned((^$unsigned(reg45)))});
          reg328 <= $signed((!{(~&reg61[(1'h1):(1'h0)]),
              $unsigned((reg18 == wire31))}));
          if ($signed($signed(reg27)))
            begin
              reg329 <= $signed(reg14[(4'hc):(3'h7)]);
            end
          else
            begin
              reg329 <= $signed($unsigned((~&$unsigned({wire324}))));
              reg330 <= $unsigned({reg20[(1'h0):(1'h0)],
                  (wire30[(4'hb):(4'hb)] < (^$signed((8'ha2))))});
              reg331 <= (!$unsigned($signed($signed((~^reg328)))));
              reg332 <= ((^$signed(((reg52 >> reg28) && {(8'ha6),
                  reg43}))) <= $signed(reg60[(4'h9):(3'h7)]));
              reg333 <= reg59[(1'h0):(1'h0)];
            end
          reg334 <= {$unsigned((wire197[(3'h7):(1'h0)] ?
                  ($unsigned(reg57) ?
                      $unsigned(reg330) : reg331) : {(reg7 && reg330),
                      reg39[(3'h7):(3'h6)]})),
              wire34};
        end
      else
        begin
          reg327 <= (wire5 ?
              $unsigned(($unsigned((wire1 ? reg14 : reg18)) ?
                  ((8'had) | reg60[(2'h2):(1'h1)]) : (^(&reg13)))) : $unsigned(($signed($unsigned(reg37)) ?
                  reg55 : reg15[(4'h8):(3'h6)])));
          reg328 <= ((wire30[(3'h6):(2'h3)] ?
                  reg8[(4'ha):(4'ha)] : reg27[(4'hd):(4'h9)]) ?
              wire2[(5'h12):(3'h6)] : (~|reg55));
          reg329 <= (reg51[(2'h3):(2'h3)] ?
              $signed((reg12[(2'h3):(1'h0)] != (reg36 ?
                  {reg39} : (reg45 > reg17)))) : (reg328 ?
                  (8'hbc) : (+$unsigned(wire4[(1'h1):(1'h1)]))));
        end
      reg335 <= reg25[(2'h3):(2'h2)];
      reg336 <= {(wire1[(1'h1):(1'h1)] ?
              ({reg331[(1'h0):(1'h0)]} ?
                  (8'hb0) : (reg21 ?
                      $signed(wire35) : (|reg16))) : (&(^~$signed((8'ha6))))),
          reg55};
      reg337 <= ((($signed($signed(wire2)) ?
          reg59[(3'h6):(1'h1)] : (((8'hb6) ? reg12 : reg9) ?
              (wire6 > reg335) : (~&reg25))) * (reg333[(4'hf):(4'hc)] ?
          ($signed(reg37) ?
              $unsigned(wire30) : (~|wire32)) : {reg18[(1'h1):(1'h1)],
              (~|wire34)})) && wire32[(2'h2):(1'h1)]);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module198
#( parameter param322 = ((({((8'h9e) >= (8'ha1))} ? (((8'ha7) ? (8'hb6) : (8'haa)) <= (+(8'hbb))) : (&{(8'ha1), (8'hb1)})) ? ((((8'hbc) ? (8'hb7) : (8'hbb)) ? {(8'hb9), (8'ha2)} : ((8'ha7) ? (8'had) : (8'ha9))) ? {((8'hb0) && (8'hbd)), (-(8'hab))} : (((8'hb5) <= (8'hbc)) ? {(8'haf)} : (~|(7'h42)))) : (({(7'h42)} ? (|(8'hbb)) : (8'hb9)) ? (((8'hb7) ? (8'h9e) : (8'hae)) == {(8'hbb)}) : (((8'hac) ~^ (8'hb9)) ? ((7'h43) ? (8'hbc) : (8'hbe)) : ((8'hb1) && (8'h9e))))) > ((((~(7'h44)) != ((8'h9f) + (8'hbf))) ^~ (!(!(8'h9f)))) > ({((8'hac) ? (8'hb3) : (8'had)), (-(8'hbb))} ? ((^~(8'ha0)) << (|(8'hb7))) : (|(7'h42)))))
, parameter param323 = (param322 ^ ((^(!{param322})) <<< (((param322 ? param322 : (8'hb7)) && (param322 << (8'hb0))) <<< param322))) )
(y, clk, wire199, wire200, wire201, wire202);
  output wire [(32'h1b1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire199;
  input wire [(4'ha):(1'h0)] wire200;
  input wire [(5'h11):(1'h0)] wire201;
  input wire signed [(4'ha):(1'h0)] wire202;
  wire [(3'h4):(1'h0)] wire226;
  reg signed [(4'h8):(1'h0)] reg228 = (1'h0);
  reg [(5'h15):(1'h0)] reg229 = (1'h0);
  reg [(4'h9):(1'h0)] reg230 = (1'h0);
  reg [(5'h15):(1'h0)] reg231 = (1'h0);
  reg [(5'h15):(1'h0)] reg232 = (1'h0);
  reg [(4'ha):(1'h0)] reg233 = (1'h0);
  reg [(5'h12):(1'h0)] reg234 = (1'h0);
  reg [(2'h3):(1'h0)] reg235 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg236 = (1'h0);
  reg [(5'h15):(1'h0)] reg237 = (1'h0);
  reg [(5'h11):(1'h0)] reg238 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg239 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg240 = (1'h0);
  reg [(5'h14):(1'h0)] reg241 = (1'h0);
  reg [(5'h10):(1'h0)] reg242 = (1'h0);
  reg [(4'he):(1'h0)] reg243 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg244 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg245 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg246 = (1'h0);
  reg [(5'h13):(1'h0)] reg247 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg248 = (1'h0);
  reg [(4'hd):(1'h0)] reg249 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire250;
  wire signed [(5'h14):(1'h0)] wire251;
  wire signed [(4'hd):(1'h0)] wire268;
  wire [(4'h9):(1'h0)] wire270;
  wire [(5'h13):(1'h0)] wire271;
  wire [(3'h5):(1'h0)] wire272;
  wire [(4'he):(1'h0)] wire296;
  wire [(4'ha):(1'h0)] wire298;
  wire signed [(3'h4):(1'h0)] wire299;
  wire [(4'hc):(1'h0)] wire300;
  wire [(5'h11):(1'h0)] wire301;
  wire signed [(4'hb):(1'h0)] wire320;
  assign y = {wire226,
                 reg228,
                 reg229,
                 reg230,
                 reg231,
                 reg232,
                 reg233,
                 reg234,
                 reg235,
                 reg236,
                 reg237,
                 reg238,
                 reg239,
                 reg240,
                 reg241,
                 reg242,
                 reg243,
                 reg244,
                 reg245,
                 reg246,
                 reg247,
                 reg248,
                 reg249,
                 wire250,
                 wire251,
                 wire268,
                 wire270,
                 wire271,
                 wire272,
                 wire296,
                 wire298,
                 wire299,
                 wire300,
                 wire301,
                 wire320,
                 (1'h0)};
  module203 modinst227 (wire226, clk, wire200, wire202, wire199, wire201, (8'hbc));
  always
    @(posedge clk) begin
      reg228 <= $signed({(-wire201[(4'hf):(3'h4)])});
      if ($unsigned($unsigned($signed($signed(((8'h9f) & wire200))))))
        begin
          reg229 <= $unsigned({(((wire202 >>> wire199) ?
                      (reg228 ? (8'ha0) : (8'hab)) : (^~wire200)) ?
                  $unsigned($signed(wire202)) : $unsigned(wire200[(2'h3):(2'h2)]))});
          reg230 <= $unsigned(((wire201 ?
              (wire226[(2'h3):(1'h1)] >= $signed(wire199)) : {((8'hb6) | reg229)}) >= ($unsigned($unsigned(wire226)) ?
              $unsigned($signed(wire199)) : wire199[(4'hb):(4'h8)])));
          reg231 <= $signed((&$unsigned(wire200[(2'h3):(2'h2)])));
          reg232 <= $signed(reg231[(4'he):(4'ha)]);
        end
      else
        begin
          if (($unsigned(wire202) * $unsigned(reg231[(4'h8):(1'h1)])))
            begin
              reg229 <= wire200;
              reg230 <= {reg229};
              reg231 <= reg232[(4'he):(4'hb)];
              reg232 <= (($unsigned({{reg229, wire202},
                      (wire226 ? wire199 : wire202)}) ?
                  (|wire226[(2'h3):(1'h0)]) : reg232) - $signed($signed(wire202[(4'ha):(2'h3)])));
              reg233 <= $signed($unsigned((~&(8'hb1))));
            end
          else
            begin
              reg229 <= $unsigned(wire200);
            end
          reg234 <= $unsigned($signed((~&$signed($unsigned(wire226)))));
          if (wire199)
            begin
              reg235 <= reg231[(5'h13):(3'h6)];
              reg236 <= $unsigned((($unsigned((reg235 ? reg231 : wire200)) ?
                      reg228 : $unsigned((~reg229))) ?
                  $signed(((~reg229) ^ $signed((8'hb0)))) : ((wire199 >>> $unsigned((8'ha2))) * {(^~wire199),
                      {wire202, reg229}})));
              reg237 <= $unsigned($signed(wire200));
            end
          else
            begin
              reg235 <= $signed({((8'ha1) ?
                      (reg235[(1'h0):(1'h0)] ?
                          wire201 : (~^reg232)) : $unsigned((wire200 ?
                          reg232 : wire202))),
                  (reg231[(4'hf):(3'h7)] >> $signed((wire226 & wire202)))});
              reg236 <= {{reg232}};
              reg237 <= (|reg237[(1'h1):(1'h0)]);
            end
          reg238 <= $unsigned(($unsigned(reg231) >> (8'ha8)));
        end
      reg239 <= reg229;
      if ((reg235[(2'h3):(2'h3)] ?
          ($signed((+$unsigned(reg228))) ?
              wire200[(3'h6):(3'h5)] : (^(~^reg232))) : (~^({(reg235 ?
                  wire200 : (8'hbb))} & ((^~wire226) ?
              (reg235 ? reg232 : (8'h9e)) : {reg235, reg233})))))
        begin
          reg240 <= $signed(reg230[(3'h6):(1'h0)]);
          if ($signed((^~{reg230[(3'h7):(3'h5)]})))
            begin
              reg241 <= (($signed(reg239[(3'h5):(1'h0)]) ?
                      wire202 : {(7'h41), reg228[(3'h7):(3'h7)]}) ?
                  (reg236 <<< $signed(wire201[(5'h10):(5'h10)])) : reg238[(4'h8):(1'h0)]);
              reg242 <= $signed((7'h43));
              reg243 <= {{(($unsigned(reg241) ?
                              $signed(reg228) : (wire226 ^ (8'hbf))) ?
                          (~&(~^wire200)) : ($unsigned(wire202) != (!reg233))),
                      $unsigned($signed($signed((8'hab))))}};
            end
          else
            begin
              reg241 <= (reg242 ?
                  $unsigned(($signed($signed((8'h9d))) >>> {(wire202 * reg228)})) : reg243[(2'h2):(2'h2)]);
              reg242 <= $signed((~(reg237 || ($signed(reg238) ?
                  ((8'hb1) ? (8'hb7) : reg233) : (~|wire226)))));
            end
          if ($signed($signed(reg238)))
            begin
              reg244 <= ((reg230[(4'h9):(1'h0)] ?
                  (~&{reg238[(2'h3):(1'h1)]}) : (-(!(reg232 >= wire199)))) >>> {({$signed(reg228)} ?
                      (~|{(8'h9d)}) : $signed((wire199 ? reg236 : reg242)))});
              reg245 <= $signed(((!(!reg241)) ?
                  {wire200, ((reg240 + reg244) << (8'hb1))} : wire200));
              reg246 <= ((wire199[(1'h0):(1'h0)] | (^~wire226)) ?
                  reg230 : $signed(reg230));
            end
          else
            begin
              reg244 <= (~$signed($signed((wire226 ?
                  (wire200 ? reg237 : wire199) : (wire226 ?
                      reg243 : reg237)))));
            end
          reg247 <= $unsigned($signed($signed($signed($unsigned(reg230)))));
        end
      else
        begin
          if ((8'hb7))
            begin
              reg240 <= {wire202[(1'h0):(1'h0)]};
              reg241 <= $unsigned((($signed($signed((8'hb0))) ?
                      ($signed(wire199) < (reg234 | reg236)) : reg233[(2'h2):(1'h0)]) ?
                  ((reg237[(4'h8):(3'h4)] ? (8'hb5) : wire200) ?
                      $signed(reg235[(2'h3):(2'h3)]) : wire226[(2'h3):(1'h1)]) : (-{$unsigned(reg243)})));
              reg242 <= ((8'haf) ?
                  (|($signed(reg247[(4'h9):(4'h9)]) ?
                      (^~((8'ha8) != reg243)) : (~(wire199 >= wire200)))) : $signed((~wire201[(4'hc):(1'h0)])));
              reg243 <= ({{($signed(wire202) + (reg232 >= reg244)),
                      reg247}} - (wire200[(1'h1):(1'h0)] | reg231[(3'h7):(1'h1)]));
              reg244 <= $unsigned((($unsigned((reg235 ? reg241 : reg242)) ?
                      $signed((reg229 | reg235)) : {reg229[(4'ha):(2'h2)]}) ?
                  $unsigned($unsigned((reg244 && (8'ha3)))) : $signed((-(~|reg229)))));
            end
          else
            begin
              reg240 <= (^(reg238 ? (-$unsigned($unsigned(reg245))) : (8'hb1)));
              reg241 <= wire199;
              reg242 <= wire202[(4'ha):(3'h7)];
            end
          if (reg247[(4'hb):(4'ha)])
            begin
              reg245 <= reg234;
              reg246 <= ($unsigned($signed($signed(reg245))) ?
                  reg244[(1'h0):(1'h0)] : (reg242 ?
                      reg235 : ($signed((reg245 ?
                          reg240 : reg244)) == $signed(reg230[(3'h7):(1'h0)]))));
            end
          else
            begin
              reg245 <= $signed(reg243);
              reg246 <= (reg239 ?
                  (reg231 <<< {$unsigned((reg245 || (8'had))),
                      ((reg245 + wire199) | (reg232 ?
                          reg244 : reg236))}) : (~&({reg245[(2'h2):(1'h0)],
                          $unsigned(reg239)} ?
                      (~&wire200[(3'h6):(3'h6)]) : ((8'h9f) ^ (reg246 ?
                          wire201 : reg243)))));
            end
          reg247 <= $signed($unsigned($unsigned((&$signed((8'hb8))))));
          reg248 <= $signed((~reg239[(3'h5):(2'h3)]));
          reg249 <= {$unsigned(reg248)};
        end
    end
  assign wire250 = {((~&($unsigned(reg249) ^~ (reg233 <= reg249))) ?
                           (~^$unsigned(reg245[(3'h5):(1'h0)])) : $signed($signed($unsigned(reg245))))};
  assign wire251 = (reg233[(3'h6):(2'h3)] ?
                       (~&($unsigned(reg241[(4'h8):(2'h3)]) && (|((8'hac) * (8'hb6))))) : (~($unsigned({reg248}) < reg237)));
  module252 modinst269 (.wire253(reg232), .clk(clk), .wire254(reg249), .wire256(wire200), .y(wire268), .wire255(reg229));
  assign wire270 = (reg233 ^~ (~^$unsigned((reg245[(2'h2):(2'h2)] >>> $unsigned(reg238)))));
  assign wire271 = (!((((reg238 * wire199) ?
                               reg235[(1'h1):(1'h1)] : (wire199 ?
                                   reg238 : reg232)) ?
                           ((-reg232) ?
                               (reg237 && reg242) : (wire251 <= wire251)) : ($signed((8'hb2)) + $unsigned(reg244))) ?
                       {wire268} : ((~^(7'h44)) >>> $signed((reg246 ?
                           (8'hb2) : reg239)))));
  assign wire272 = ($signed((((reg235 ? wire250 : reg231) ?
                               $signed(reg241) : (reg249 >>> reg245)) ?
                           (~^$unsigned(reg240)) : (reg228[(3'h6):(2'h2)] | $unsigned((8'hba))))) ?
                       reg249[(4'hb):(3'h5)] : {$unsigned(((reg247 ~^ wire250) ?
                               $signed((8'ha7)) : $unsigned(reg249)))});
  module273 modinst297 (.wire276(reg242), .wire277(wire202), .wire274(wire251), .y(wire296), .wire275(reg243), .clk(clk));
  assign wire298 = ($unsigned(((8'hb1) <= $signed($unsigned((7'h41))))) < $signed($signed({(wire199 ?
                           reg245 : reg248),
                       $signed(wire199)})));
  assign wire299 = reg238[(3'h5):(3'h5)];
  assign wire300 = reg237;
  assign wire301 = {reg248};
  module302 modinst321 (wire320, clk, reg232, wire298, reg237, reg238, reg248);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module66
#( parameter param194 = ((((((7'h41) ? (8'h9d) : (8'hb3)) || (&(8'h9f))) ? (~&((8'hba) <<< (8'ha8))) : (((8'ha2) < (7'h40)) | ((8'hbb) == (8'hb7)))) << (+(((8'ha8) ? (8'ha7) : (8'hac)) && (8'ha9)))) ~^ {({(~^(8'h9c)), ((7'h41) ^ (8'hbd))} ? (((8'ha4) ? (8'hbc) : (8'hab)) < ((8'hb7) ^ (8'haf))) : (^(8'hab)))}) )
(y, clk, wire67, wire68, wire69, wire70, wire71);
  output wire [(32'h135):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire67;
  input wire [(4'hd):(1'h0)] wire68;
  input wire signed [(4'h9):(1'h0)] wire69;
  input wire [(3'h7):(1'h0)] wire70;
  input wire signed [(4'hf):(1'h0)] wire71;
  wire signed [(4'hd):(1'h0)] wire193;
  wire signed [(4'hf):(1'h0)] wire72;
  wire [(5'h15):(1'h0)] wire73;
  wire signed [(4'hf):(1'h0)] wire74;
  wire signed [(4'he):(1'h0)] wire75;
  wire [(4'hc):(1'h0)] wire76;
  wire signed [(4'h9):(1'h0)] wire77;
  wire signed [(4'he):(1'h0)] wire78;
  wire [(5'h12):(1'h0)] wire79;
  wire signed [(5'h13):(1'h0)] wire80;
  reg signed [(5'h13):(1'h0)] reg81 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg82 = (1'h0);
  reg [(3'h4):(1'h0)] reg83 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg84 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg85 = (1'h0);
  reg [(4'hd):(1'h0)] reg86 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg87 = (1'h0);
  wire [(3'h7):(1'h0)] wire88;
  reg signed [(3'h6):(1'h0)] reg89 = (1'h0);
  reg [(3'h6):(1'h0)] reg90 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire91;
  wire signed [(4'h8):(1'h0)] wire111;
  wire signed [(4'hc):(1'h0)] wire113;
  wire signed [(4'hd):(1'h0)] wire114;
  wire [(5'h11):(1'h0)] wire191;
  assign y = {wire193,
                 wire72,
                 wire73,
                 wire74,
                 wire75,
                 wire76,
                 wire77,
                 wire78,
                 wire79,
                 wire80,
                 reg81,
                 reg82,
                 reg83,
                 reg84,
                 reg85,
                 reg86,
                 reg87,
                 wire88,
                 reg89,
                 reg90,
                 wire91,
                 wire111,
                 wire113,
                 wire114,
                 wire191,
                 (1'h0)};
  assign wire72 = wire67[(5'h14):(4'h8)];
  assign wire73 = $signed((~^($unsigned($unsigned(wire68)) || ($signed(wire68) < (~|wire67)))));
  assign wire74 = $unsigned(wire68);
  assign wire75 = wire69;
  assign wire76 = wire69[(4'h9):(1'h0)];
  assign wire77 = $unsigned(($signed($unsigned(wire70[(2'h2):(1'h0)])) & wire67[(3'h6):(3'h6)]));
  assign wire78 = (&$signed(((!(~|wire69)) ? wire77 : wire73[(4'hd):(3'h4)])));
  assign wire79 = $signed($signed(({wire75} ? wire68 : {$unsigned(wire67)})));
  assign wire80 = wire70;
  always
    @(posedge clk) begin
      if (((wire67 >> wire77[(4'h9):(2'h2)]) >> $unsigned((!$unsigned(((8'ha9) ?
          (8'h9d) : wire80))))))
        begin
          reg81 <= (|($signed((wire77[(2'h3):(1'h0)] >>> wire68)) + ((wire74[(4'ha):(1'h0)] ?
                  wire73[(5'h11):(2'h3)] : $signed(wire70)) ?
              $signed($unsigned(wire79)) : wire71[(4'hf):(4'hc)])));
        end
      else
        begin
          reg81 <= $signed(wire75[(4'ha):(4'h8)]);
          reg82 <= (wire78[(1'h0):(1'h0)] ?
              $signed(wire78) : ($signed((^~(!wire76))) ?
                  $signed(($unsigned(wire70) || (wire75 || wire71))) : ($unsigned($signed(wire79)) ?
                      (-wire71[(4'hd):(4'hb)]) : ({wire74,
                          wire80} - (wire77 ^~ wire67)))));
        end
      if (reg82[(1'h0):(1'h0)])
        begin
          reg83 <= ({(&((!reg82) <= (wire79 ? wire70 : wire79))),
              wire80[(4'hd):(1'h1)]} <= ((8'hb9) ?
              (+wire77[(3'h5):(2'h3)]) : $unsigned(({wire79} ?
                  (wire75 | (8'hae)) : $signed(wire72)))));
          reg84 <= (wire70[(3'h4):(1'h1)] & {{((wire78 - wire67) ?
                      (wire67 || (8'hb2)) : wire70)}});
          reg85 <= ($signed(($unsigned((wire70 ? wire78 : wire79)) ?
                  wire75 : (~wire69[(4'h9):(1'h0)]))) ?
              $signed((wire76[(2'h2):(2'h2)] >> $signed((~^(8'ha7))))) : (+wire77));
          reg86 <= (-$unsigned(($signed((reg83 ?
              reg83 : wire75)) ~^ ((&(8'hb8)) ? reg83 : (|wire74)))));
        end
      else
        begin
          reg83 <= $unsigned($signed(wire67[(5'h11):(4'hc)]));
        end
      reg87 <= wire71;
    end
  assign wire88 = wire74[(4'h9):(2'h3)];
  always
    @(posedge clk) begin
      reg89 <= wire70[(2'h3):(2'h2)];
      reg90 <= wire70;
    end
  assign wire91 = reg89[(2'h2):(1'h1)];
  module92 modinst112 (.wire93(wire72), .wire94(reg81), .wire95(wire88), .clk(clk), .y(wire111), .wire96(wire74));
  assign wire113 = {($unsigned(($unsigned(reg87) == ((8'hb3) | wire76))) != $unsigned(((reg81 ?
                           wire68 : (8'haf)) >>> wire75[(3'h6):(2'h3)])))};
  assign wire114 = reg90[(1'h1):(1'h1)];
  module115 modinst192 (.y(wire191), .clk(clk), .wire119(wire78), .wire120(wire91), .wire117(wire68), .wire116(reg81), .wire118(wire74));
  assign wire193 = (~wire88);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module115
#( parameter param190 = ({((((8'h9e) ? (8'hbb) : (8'hac)) < (^(8'ha3))) >>> ((&(8'ha9)) ? ((8'hb8) && (8'hbc)) : (^~(8'ha1))))} - (~&((((8'h9f) << (8'h9c)) ? ((7'h44) * (8'hbf)) : (8'hac)) ^ {{(8'ha6), (8'hbc)}, ((8'hac) ? (8'hbb) : (8'hab))}))) )
(y, clk, wire120, wire119, wire118, wire117, wire116);
  output wire [(32'h332):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h6):(1'h0)] wire120;
  input wire signed [(3'h4):(1'h0)] wire119;
  input wire [(3'h5):(1'h0)] wire118;
  input wire [(4'hd):(1'h0)] wire117;
  input wire signed [(2'h2):(1'h0)] wire116;
  wire signed [(5'h12):(1'h0)] wire189;
  wire signed [(5'h11):(1'h0)] wire188;
  reg signed [(5'h15):(1'h0)] reg187 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg186 = (1'h0);
  reg [(5'h11):(1'h0)] reg185 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg184 = (1'h0);
  reg [(4'h8):(1'h0)] reg183 = (1'h0);
  reg [(3'h7):(1'h0)] reg182 = (1'h0);
  reg [(4'h9):(1'h0)] reg181 = (1'h0);
  reg [(5'h11):(1'h0)] reg180 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg179 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg178 = (1'h0);
  reg [(5'h12):(1'h0)] reg177 = (1'h0);
  reg [(5'h10):(1'h0)] reg176 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg175 = (1'h0);
  reg [(3'h5):(1'h0)] reg174 = (1'h0);
  reg [(4'ha):(1'h0)] reg173 = (1'h0);
  reg [(4'hd):(1'h0)] reg172 = (1'h0);
  reg [(3'h4):(1'h0)] reg171 = (1'h0);
  reg [(5'h11):(1'h0)] reg170 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg169 = (1'h0);
  reg [(4'hb):(1'h0)] reg168 = (1'h0);
  reg [(4'h9):(1'h0)] reg167 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg166 = (1'h0);
  reg [(5'h14):(1'h0)] reg165 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg164 = (1'h0);
  reg [(3'h4):(1'h0)] reg163 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg162 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire161;
  wire signed [(4'h9):(1'h0)] wire160;
  wire signed [(3'h7):(1'h0)] wire159;
  wire signed [(4'h8):(1'h0)] wire158;
  wire [(3'h5):(1'h0)] wire157;
  reg [(4'h9):(1'h0)] reg156 = (1'h0);
  reg [(2'h2):(1'h0)] reg155 = (1'h0);
  reg [(3'h7):(1'h0)] reg154 = (1'h0);
  reg signed [(4'he):(1'h0)] reg153 = (1'h0);
  reg [(4'hb):(1'h0)] reg152 = (1'h0);
  reg [(4'hb):(1'h0)] reg151 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg150 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg149 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg148 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg147 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg146 = (1'h0);
  reg [(4'he):(1'h0)] reg145 = (1'h0);
  reg [(4'hf):(1'h0)] reg144 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg143 = (1'h0);
  reg [(4'he):(1'h0)] reg142 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg141 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg140 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg139 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg138 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg137 = (1'h0);
  reg [(4'h8):(1'h0)] reg136 = (1'h0);
  reg [(5'h11):(1'h0)] reg135 = (1'h0);
  reg signed [(4'he):(1'h0)] reg134 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg133 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg132 = (1'h0);
  reg [(5'h11):(1'h0)] reg131 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg130 = (1'h0);
  reg [(4'h8):(1'h0)] reg129 = (1'h0);
  wire [(4'hd):(1'h0)] wire128;
  wire signed [(3'h4):(1'h0)] wire127;
  wire [(3'h4):(1'h0)] wire126;
  wire [(5'h15):(1'h0)] wire125;
  wire [(4'hc):(1'h0)] wire124;
  wire [(5'h13):(1'h0)] wire123;
  wire signed [(3'h7):(1'h0)] wire122;
  wire [(2'h3):(1'h0)] wire121;
  assign y = {wire189,
                 wire188,
                 reg187,
                 reg186,
                 reg185,
                 reg184,
                 reg183,
                 reg182,
                 reg181,
                 reg180,
                 reg179,
                 reg178,
                 reg177,
                 reg176,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 wire161,
                 wire160,
                 wire159,
                 wire158,
                 wire157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 reg149,
                 reg148,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 reg143,
                 reg142,
                 reg141,
                 reg140,
                 reg139,
                 reg138,
                 reg137,
                 reg136,
                 reg135,
                 reg134,
                 reg133,
                 reg132,
                 reg131,
                 reg130,
                 reg129,
                 wire128,
                 wire127,
                 wire126,
                 wire125,
                 wire124,
                 wire123,
                 wire122,
                 wire121,
                 (1'h0)};
  assign wire121 = wire120[(3'h6):(2'h3)];
  assign wire122 = wire121[(1'h0):(1'h0)];
  assign wire123 = wire122[(3'h5):(3'h5)];
  assign wire124 = wire119;
  assign wire125 = $unsigned(wire116);
  assign wire126 = $unsigned($signed(({wire118} ?
                       ($signed(wire118) ?
                           wire125 : $unsigned(wire123)) : wire118)));
  assign wire127 = (-(~^{wire116[(1'h1):(1'h1)],
                       (wire124[(4'hb):(4'hb)] > (wire119 ?
                           wire124 : wire118))}));
  assign wire128 = $signed({$unsigned(((wire124 ? wire126 : wire125) ?
                           wire127 : (wire127 >> (8'h9d)))),
                       wire118});
  always
    @(posedge clk) begin
      reg129 <= (~$signed((wire123[(2'h3):(2'h3)] ?
          ((wire120 + wire122) <<< $signed(wire120)) : wire121[(2'h2):(1'h1)])));
      reg130 <= (-$signed($unsigned($unsigned(((8'ha6) ? (8'hb1) : wire119)))));
      reg131 <= reg129;
      reg132 <= (8'ha4);
      if ((wire128 << reg132[(3'h6):(1'h0)]))
        begin
          reg133 <= $unsigned($unsigned(({{wire122, wire121},
                  (wire116 ^ wire119)} ?
              (reg129[(3'h4):(3'h4)] * (^(8'had))) : $signed((^(8'hbd))))));
          if ((8'ha6))
            begin
              reg134 <= ($signed(wire125[(3'h6):(3'h6)]) ?
                  (reg130[(1'h1):(1'h1)] <= (((reg130 != wire119) | (wire125 ?
                          wire128 : (8'had))) ?
                      wire125[(1'h0):(1'h0)] : $unsigned((~&wire126)))) : reg131);
              reg135 <= $unsigned(wire117[(3'h6):(3'h5)]);
              reg136 <= ((wire128[(1'h0):(1'h0)] ?
                      (((!(8'hb4)) >> reg135[(3'h4):(2'h2)]) ?
                          ((reg130 - reg135) ?
                              reg132[(3'h6):(1'h1)] : (wire122 ?
                                  reg130 : wire116)) : wire123) : $unsigned(wire118)) ?
                  (&reg129) : (reg134[(4'hb):(3'h6)] > (reg135 ?
                      {(wire123 ? wire116 : (8'hbc))} : (+(wire123 ?
                          wire124 : reg133)))));
            end
          else
            begin
              reg134 <= $unsigned(($signed((wire125 >= (wire116 * wire116))) + {wire122,
                  wire122[(1'h1):(1'h1)]}));
              reg135 <= wire118;
              reg136 <= ($unsigned(($signed((~wire117)) || $unsigned(wire123[(5'h13):(1'h0)]))) ?
                  {$signed({$signed(wire119),
                          {reg135, (8'hba)}})} : ($signed((|$signed((8'ha2)))) ?
                      $unsigned((reg136[(3'h6):(3'h5)] << (wire117 ?
                          (8'hb7) : wire119))) : $unsigned(wire127)));
              reg137 <= reg129[(3'h6):(1'h0)];
            end
          if ((!{$unsigned(({wire127} < (wire120 >>> wire118))),
              ({(!reg134)} | wire121[(1'h1):(1'h0)])}))
            begin
              reg138 <= $signed($unsigned(reg137));
              reg139 <= reg138[(3'h7):(3'h4)];
              reg140 <= reg139;
              reg141 <= ($unsigned(($signed((wire124 + reg140)) && ((reg139 <= reg132) != (!reg134)))) ?
                  reg131 : $unsigned($unsigned(((wire118 ?
                      (8'hbd) : reg132) != (8'haf)))));
              reg142 <= (((reg135 ?
                  $unsigned(wire121[(2'h3):(1'h1)]) : ($unsigned(reg140) > (reg132 ?
                      wire120 : wire119))) || wire120) || (reg132 ?
                  (reg133 || reg136) : reg140[(5'h12):(5'h11)]));
            end
          else
            begin
              reg138 <= (&wire117[(1'h0):(1'h0)]);
              reg139 <= wire119[(2'h3):(2'h2)];
              reg140 <= $unsigned(((8'hba) ? wire120 : reg131[(4'ha):(4'ha)]));
            end
        end
      else
        begin
          reg133 <= $unsigned((~|$unsigned($signed((reg134 ?
              (8'hbd) : (8'hb5))))));
        end
    end
  always
    @(posedge clk) begin
      reg143 <= wire122;
      reg144 <= (^~wire127);
      reg145 <= (!$unsigned($signed(wire128[(4'ha):(3'h6)])));
    end
  always
    @(posedge clk) begin
      reg146 <= (!$signed($unsigned((reg134 ?
          reg138[(3'h7):(2'h3)] : (!reg145)))));
      if ({$signed({wire126[(2'h3):(1'h0)]})})
        begin
          reg147 <= (((reg138 >= reg140) != reg141[(1'h1):(1'h0)]) >>> reg137);
          reg148 <= {wire126[(3'h4):(1'h0)]};
          reg149 <= wire122[(3'h5):(2'h2)];
        end
      else
        begin
          reg147 <= ($unsigned((-($signed(reg145) ?
              {reg140, reg139} : $signed(reg129)))) + (-reg141[(2'h3):(2'h2)]));
          if (reg143)
            begin
              reg148 <= wire116[(1'h1):(1'h0)];
              reg149 <= wire123[(4'h8):(3'h4)];
              reg150 <= wire125;
            end
          else
            begin
              reg148 <= ({$unsigned((+{reg129, reg134})),
                  $signed(reg148[(4'he):(2'h3)])} != $unsigned({reg145}));
              reg149 <= reg149;
              reg150 <= $unsigned(($unsigned(reg135[(4'ha):(2'h3)]) ?
                  $unsigned(reg140) : reg141[(1'h1):(1'h0)]));
              reg151 <= $signed({(^~{(reg136 ? (8'ha5) : reg136), reg140}),
                  (8'hb9)});
            end
          if ((-(~^reg142)))
            begin
              reg152 <= (-wire119[(3'h4):(2'h3)]);
              reg153 <= reg129[(3'h7):(3'h7)];
              reg154 <= reg151;
              reg155 <= ($unsigned((((&wire123) ?
                  (reg150 ?
                      wire123 : (8'h9c)) : reg144[(3'h4):(1'h0)]) ~^ $unsigned((reg141 ?
                  reg134 : reg135)))) >> (reg133[(4'hc):(1'h1)] ?
                  ($signed((reg152 ? reg147 : reg144)) ?
                      (reg141 ?
                          $unsigned(reg148) : reg139[(4'hb):(4'ha)]) : ({(8'hbf)} ^ (wire127 || wire123))) : $signed($unsigned($unsigned((8'hb5))))));
            end
          else
            begin
              reg152 <= wire117[(3'h5):(1'h1)];
              reg153 <= reg148[(5'h15):(2'h3)];
              reg154 <= ((&(+($unsigned(reg136) ?
                  $unsigned(wire121) : wire117))) + (~&((8'ha5) ?
                  wire121[(1'h0):(1'h0)] : $signed($signed(wire127)))));
              reg155 <= $unsigned(reg149[(3'h7):(1'h1)]);
            end
        end
      reg156 <= wire118[(1'h1):(1'h0)];
    end
  assign wire157 = (((((!reg144) ?
                           (reg129 ?
                               wire122 : reg137) : (reg143 || wire119)) != (reg156 ~^ wire121)) ?
                       (!(~&$unsigned((8'hbe)))) : $signed(((~|reg149) <<< reg133[(4'hb):(4'h8)]))) > ($signed($signed($unsigned(reg142))) >>> (reg131[(3'h6):(3'h4)] ?
                       {(wire123 ~^ reg145)} : (~&$signed(wire121)))));
  assign wire158 = $signed((({((7'h44) != wire157), $unsigned((8'hb0))} ?
                           (-(~&reg149)) : ((8'ha7) - reg132[(4'h8):(1'h1)])) ?
                       ((-(wire128 ? reg153 : wire122)) ?
                           (((8'h9c) ?
                               wire124 : (7'h40)) != (reg130 >>> reg138)) : {(reg135 ?
                                   reg140 : reg136),
                               reg148[(5'h15):(4'h9)]}) : $unsigned({(wire116 ?
                               wire123 : reg141)})));
  assign wire159 = {($signed(((reg129 && reg150) ^~ $signed(reg147))) && (&$signed(wire128))),
                       {(reg148[(4'hc):(4'h9)] ?
                               $signed((reg145 >= reg156)) : wire118[(2'h2):(2'h2)]),
                           (wire126[(2'h3):(2'h3)] ?
                               (^{reg136}) : $signed((8'ha6)))}};
  assign wire160 = (wire119[(2'h2):(1'h1)] << wire117[(3'h5):(2'h2)]);
  assign wire161 = $unsigned((-$signed(((reg134 * (8'hb5)) ?
                       $unsigned((8'haa)) : reg151[(4'hb):(3'h4)]))));
  always
    @(posedge clk) begin
      if ($signed($signed((~^(+$unsigned(reg131))))))
        begin
          reg162 <= $unsigned($unsigned($signed(((wire128 || (7'h43)) ?
              reg139[(1'h1):(1'h0)] : (|reg149)))));
          reg163 <= (-wire160[(3'h6):(2'h3)]);
        end
      else
        begin
          reg162 <= $signed((&$signed(reg154)));
          if ((|{(&(^~wire124[(1'h0):(1'h0)])),
              $signed($signed($signed(reg162)))}))
            begin
              reg163 <= wire157[(2'h3):(1'h0)];
              reg164 <= ((~(&wire116)) ?
                  (-wire117[(3'h5):(1'h1)]) : $signed(($unsigned({reg131,
                          (8'hbd)}) ?
                      $unsigned({reg142, wire125}) : reg149[(4'h8):(1'h0)])));
              reg165 <= (((!((wire117 >>> (8'hbf)) ?
                  wire157 : (^~reg163))) <<< ($unsigned($signed((7'h43))) ?
                  reg138[(1'h1):(1'h0)] : reg151[(4'h8):(3'h4)])) + (reg164 || reg164));
              reg166 <= (wire124 ? wire118[(1'h0):(1'h0)] : wire126);
              reg167 <= (($unsigned(wire123[(3'h5):(2'h2)]) && $unsigned(((reg142 ?
                      reg135 : wire127) ?
                  $signed(reg129) : wire125))) <= (^~($unsigned({reg140,
                  wire122}) ~^ $signed((wire121 - reg139)))));
            end
          else
            begin
              reg163 <= ($unsigned($unsigned(((8'ha0) ?
                  {(8'ha4), reg143} : (reg136 ?
                      (8'hb3) : (8'hba))))) ^ ($unsigned((&$unsigned(reg150))) && (^~(8'ha0))));
              reg164 <= reg156;
              reg165 <= ((reg133 ?
                  ((wire125 ? ((7'h44) ? reg135 : wire118) : wire159) ?
                      (8'hb1) : (8'hb7)) : reg145[(3'h4):(2'h3)]) >= (($signed(reg130) ?
                  wire158[(1'h1):(1'h1)] : {(8'hb7)}) | ((~$unsigned(reg163)) ?
                  (|{reg148}) : (~^(~^reg139)))));
              reg166 <= ({wire120[(3'h5):(1'h1)]} == (+((wire157[(3'h4):(1'h0)] >>> {reg166,
                  (8'haf)}) * reg140[(1'h0):(1'h0)])));
            end
          reg168 <= {reg141, (|{($signed(reg145) * reg145)})};
          reg169 <= ($unsigned(((8'h9f) ?
                  wire128 : (~|reg155[(1'h1):(1'h1)]))) ?
              (|(reg149[(2'h3):(1'h1)] ?
                  wire157 : ((~^(8'h9d)) & $signed(reg144)))) : $unsigned((8'hbf)));
        end
    end
  always
    @(posedge clk) begin
      if ($unsigned($signed((reg151[(2'h3):(1'h0)] ?
          (~&$signed(reg142)) : ($unsigned(reg138) ?
              (reg163 * wire127) : reg163[(2'h3):(2'h2)])))))
        begin
          reg170 <= {reg167};
          reg171 <= (((8'haf) ~^ (8'had)) <= (^wire116[(1'h0):(1'h0)]));
          if ((~^(^~reg162)))
            begin
              reg172 <= $signed(($signed(wire121[(1'h1):(1'h1)]) ^ ((reg133[(3'h4):(3'h4)] ?
                  {wire120, (7'h40)} : $signed((8'ha7))) <= ((reg138 ?
                  reg156 : reg169) << (reg144 ? reg146 : reg163)))));
            end
          else
            begin
              reg172 <= $unsigned(((-((&wire120) ?
                  (reg141 ?
                      reg146 : reg151) : reg172)) != ($signed($unsigned(wire125)) ?
                  ((~&reg129) * $unsigned(wire127)) : (+{(8'hb4)}))));
              reg173 <= reg154;
              reg174 <= (^~(reg142[(4'ha):(4'ha)] ?
                  $signed(((reg130 <<< reg169) * $signed(reg130))) : ((&(reg171 < reg168)) || ($signed(reg132) ?
                      (~&reg144) : wire126[(2'h3):(1'h0)]))));
            end
        end
      else
        begin
          reg170 <= (^~reg152[(3'h5):(3'h5)]);
          reg171 <= $unsigned((~^{reg149,
              (reg173[(2'h3):(2'h2)] ?
                  reg148[(5'h12):(4'h8)] : reg172[(3'h5):(1'h1)])}));
          reg172 <= (reg169 ?
              (wire128[(2'h2):(1'h0)] ?
                  $signed({wire127}) : (^~$unsigned(((8'hbc) >>> wire125)))) : (~^(($unsigned(reg136) || ((8'hac) ~^ reg173)) | reg152[(4'h9):(3'h6)])));
        end
      reg175 <= (!$signed($signed(($unsigned(reg155) >> (-reg154)))));
      reg176 <= ((~|(+{{reg154, reg139}, $signed(reg156)})) ?
          ({(^$unsigned(wire158)),
              reg169[(3'h5):(3'h4)]} || {$unsigned(wire121[(2'h3):(2'h2)]),
              $unsigned({(8'hac)})}) : $unsigned((8'hb1)));
      reg177 <= ((~^((reg130[(1'h0):(1'h0)] <= (reg138 || reg132)) ?
          $unsigned((8'h9d)) : $signed((8'h9c)))) >= (~|($signed($unsigned(reg146)) ?
          (wire121[(1'h0):(1'h0)] ^ reg135) : (reg136[(1'h0):(1'h0)] >> (reg132 ?
              (8'hbb) : wire158)))));
      if ($unsigned((reg177[(2'h3):(1'h1)] ^ $signed($signed(reg139[(4'hf):(1'h1)])))))
        begin
          reg178 <= {$signed(reg167)};
          if ({$signed(reg147[(2'h2):(2'h2)]), (8'hba)})
            begin
              reg179 <= (~|{$signed((reg155[(1'h1):(1'h1)] < reg132[(5'h11):(5'h11)]))});
              reg180 <= ($unsigned(((~|wire158) ?
                  {(reg145 ^ (8'hb4))} : wire127)) >>> {reg134});
              reg181 <= $unsigned($signed({reg177}));
              reg182 <= ((+$unsigned(($unsigned(wire116) ?
                      (reg170 ? reg136 : wire116) : (reg162 != reg170)))) ?
                  wire128[(4'hd):(4'hd)] : (7'h44));
              reg183 <= ((~|$signed(reg132[(1'h0):(1'h0)])) ?
                  reg182 : ($unsigned($unsigned({wire161})) <<< wire126[(2'h3):(1'h0)]));
            end
          else
            begin
              reg179 <= ($unsigned((((8'h9f) * $signed(reg136)) ?
                  (~&(wire159 ?
                      reg176 : wire128)) : $unsigned($signed(reg175)))) ^ $signed($unsigned(reg139)));
              reg180 <= reg148[(3'h7):(3'h7)];
              reg181 <= $unsigned(({reg183} ^~ $signed(((reg153 ?
                      reg149 : reg131) ?
                  (reg181 ? reg171 : wire120) : $signed(reg178)))));
              reg182 <= (&reg154[(3'h4):(2'h3)]);
            end
          if ((~&$unsigned($unsigned(((reg143 ? wire117 : reg166) ?
              $signed((8'had)) : $signed((8'had)))))))
            begin
              reg184 <= (^~((($signed(wire128) ?
                          (wire118 ? reg167 : (8'hbf)) : (wire119 ?
                              reg180 : reg151)) ?
                      reg141[(1'h1):(1'h0)] : reg142[(4'h9):(3'h6)]) ?
                  ((~^(~&wire120)) >> $unsigned((~wire118))) : reg132[(3'h6):(2'h2)]));
              reg185 <= (wire128[(4'hd):(2'h2)] ?
                  ($signed(($unsigned(reg184) ?
                      (wire161 ?
                          reg133 : (8'haa)) : $signed(reg177))) != ({$unsigned(reg142),
                          $unsigned(reg150)} ?
                      ((reg143 == wire120) ?
                          ((8'hb1) ?
                              (8'h9d) : wire124) : (reg133 != reg155)) : reg133)) : reg162);
              reg186 <= $signed(($signed((wire122 ?
                      $signed(reg179) : {reg129})) ?
                  ($signed(wire121) ?
                      $unsigned((8'ha7)) : ((reg177 >> reg147) ?
                          $signed((8'hb3)) : (reg177 | reg145))) : (^(-(wire116 ?
                      wire124 : reg147)))));
            end
          else
            begin
              reg184 <= (((((reg143 * reg150) * reg171) != ((reg150 ?
                              reg186 : wire118) ?
                          (wire120 ^ reg155) : (reg176 ? reg156 : (7'h41)))) ?
                      (reg162 ?
                          (8'hac) : ($signed((8'hb7)) ?
                              $unsigned(reg185) : reg145)) : (~(reg181 ?
                          reg165 : (|wire117)))) ?
                  $unsigned(((wire125 ? reg154 : reg171[(2'h3):(1'h0)]) ?
                      {(reg185 ?
                              reg165 : reg176)} : (reg167[(4'h9):(4'h8)] & $signed((8'h9f))))) : $signed((reg142 <<< $signed((^~reg141)))));
            end
          reg187 <= reg150;
        end
      else
        begin
          reg178 <= $unsigned($unsigned(($unsigned(reg147[(1'h0):(1'h0)]) ?
              reg156 : reg144[(3'h5):(1'h0)])));
          if (reg173)
            begin
              reg179 <= (($signed(($signed(reg147) ?
                          $unsigned((8'hab)) : reg135)) ?
                      $unsigned(($signed((8'h9f)) & (wire120 ?
                          wire123 : reg140))) : (~(&$signed(reg151)))) ?
                  (+reg130) : $unsigned($unsigned($signed((reg142 ~^ wire158)))));
              reg180 <= {reg180};
            end
          else
            begin
              reg179 <= reg155[(1'h1):(1'h1)];
              reg180 <= (!(reg170 ?
                  (~((reg175 ? (8'hb4) : reg133) <= (~wire122))) : reg131));
              reg181 <= ($signed($unsigned(((reg170 << (8'hb0)) & (reg162 == reg186)))) & {reg154,
                  (reg184[(2'h2):(1'h0)] ?
                      (+reg142[(4'h9):(3'h7)]) : (-(+reg141)))});
              reg182 <= (!{$unsigned(reg162[(4'h9):(3'h6)])});
            end
          reg183 <= (&wire120);
          reg184 <= ($unsigned((((reg137 <<< reg131) & $unsigned(reg174)) | reg145)) == $signed(reg167));
        end
    end
  assign wire188 = $unsigned({(($signed(reg177) <= $unsigned((8'ha2))) ?
                           $signed($unsigned(reg184)) : reg182[(3'h6):(2'h2)]),
                       reg141});
  assign wire189 = (($unsigned((|(-wire117))) ?
                       ({((7'h42) ? wire119 : reg180),
                           (!reg173)} ^ ($signed(reg143) || (reg155 << (8'h9e)))) : (wire188 + $signed((reg187 ^~ reg154)))) ^ $unsigned(($unsigned(reg167) ?
                       $signed(wire125[(5'h11):(1'h1)]) : ((reg140 + reg168) >>> $unsigned(reg148)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module92
#( parameter param110 = {(~&(~&({(8'ha6)} ? ((8'ha7) ? (8'hba) : (8'hbd)) : {(8'haf), (8'ha2)})))} )
(y, clk, wire96, wire95, wire94, wire93);
  output wire [(32'h80):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h5):(1'h0)] wire96;
  input wire [(2'h3):(1'h0)] wire95;
  input wire [(5'h13):(1'h0)] wire94;
  input wire signed [(4'h8):(1'h0)] wire93;
  wire [(2'h2):(1'h0)] wire109;
  wire [(3'h5):(1'h0)] wire108;
  wire signed [(4'hf):(1'h0)] wire107;
  reg [(4'ha):(1'h0)] reg106 = (1'h0);
  reg [(4'h9):(1'h0)] reg105 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg104 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire103;
  wire [(3'h6):(1'h0)] wire102;
  wire signed [(4'ha):(1'h0)] wire101;
  wire signed [(4'ha):(1'h0)] wire100;
  wire signed [(2'h3):(1'h0)] wire99;
  wire signed [(5'h14):(1'h0)] wire98;
  wire [(5'h14):(1'h0)] wire97;
  assign y = {wire109,
                 wire108,
                 wire107,
                 reg106,
                 reg105,
                 reg104,
                 wire103,
                 wire102,
                 wire101,
                 wire100,
                 wire99,
                 wire98,
                 wire97,
                 (1'h0)};
  assign wire97 = $signed(wire96[(3'h5):(1'h1)]);
  assign wire98 = ((wire96[(2'h3):(1'h0)] ~^ wire95) ?
                      $unsigned((8'hb7)) : ((^{wire95[(1'h0):(1'h0)], wire97}) ?
                          (!$unsigned(wire97)) : ($unsigned(wire95) ?
                              ($signed(wire94) ?
                                  (wire95 ?
                                      wire95 : wire93) : (+wire96)) : wire97)));
  assign wire99 = wire98[(1'h0):(1'h0)];
  assign wire100 = wire99[(2'h2):(1'h0)];
  assign wire101 = $unsigned(wire96[(3'h5):(2'h3)]);
  assign wire102 = $unsigned(wire101[(4'ha):(3'h4)]);
  assign wire103 = (((8'h9c) == $signed(wire96[(2'h2):(1'h0)])) ?
                       $signed((~^($signed(wire100) || (wire101 <= wire95)))) : ($signed(((^wire98) ?
                               (^wire99) : (|wire95))) ?
                           wire93 : $unsigned(wire94)));
  always
    @(posedge clk) begin
      reg104 <= {{wire93}, wire99};
      reg105 <= wire97[(4'hb):(3'h5)];
      reg106 <= $unsigned({wire100});
    end
  assign wire107 = $unsigned(({wire101, (~|wire103)} ?
                       $signed(((^~reg105) ?
                           reg106[(4'h9):(1'h0)] : wire96[(1'h0):(1'h0)])) : reg104));
  assign wire108 = (((|$signed((wire93 ?
                       wire103 : (8'ha2)))) + wire107) | (^~$unsigned(wire96)));
  assign wire109 = wire108;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module302
#( parameter param319 = (({((^~(8'ha2)) | {(8'ha8), (8'hb0)})} ? {(((8'ha4) - (8'hb1)) ^~ ((8'hba) ^~ (8'ha8)))} : {{{(8'haa), (8'hb4)}}}) == (((7'h42) ? ((~^(8'ha4)) || (~|(8'ha2))) : (((8'hac) ? (8'hbc) : (7'h44)) ? ((8'ha1) + (8'hae)) : ((8'hbf) << (8'hb6)))) ? (8'ha7) : ((~|((7'h44) & (8'hb2))) ? ((~^(8'hb5)) != ((8'hb9) << (8'hba))) : (!((8'hae) ? (8'ha6) : (8'ha0)))))) )
(y, clk, wire307, wire306, wire305, wire304, wire303);
  output wire [(32'h86):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire307;
  input wire [(4'h9):(1'h0)] wire306;
  input wire signed [(2'h2):(1'h0)] wire305;
  input wire [(5'h11):(1'h0)] wire304;
  input wire [(2'h3):(1'h0)] wire303;
  wire [(5'h13):(1'h0)] wire318;
  wire [(5'h14):(1'h0)] wire317;
  wire [(4'ha):(1'h0)] wire316;
  wire [(5'h11):(1'h0)] wire315;
  wire signed [(2'h2):(1'h0)] wire314;
  reg signed [(4'hb):(1'h0)] reg313 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg312 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg311 = (1'h0);
  wire [(4'hd):(1'h0)] wire310;
  wire [(3'h4):(1'h0)] wire309;
  wire [(4'he):(1'h0)] wire308;
  assign y = {wire318,
                 wire317,
                 wire316,
                 wire315,
                 wire314,
                 reg313,
                 reg312,
                 reg311,
                 wire310,
                 wire309,
                 wire308,
                 (1'h0)};
  assign wire308 = (wire306[(1'h0):(1'h0)] ?
                       $signed(wire303[(2'h2):(1'h0)]) : $unsigned((-wire303[(2'h3):(1'h0)])));
  assign wire309 = wire304[(4'ha):(3'h7)];
  assign wire310 = $signed($signed($signed($unsigned(wire304))));
  always
    @(posedge clk) begin
      reg311 <= {wire309};
      reg312 <= $unsigned(wire309);
      reg313 <= (wire303 ? wire308 : (8'h9e));
    end
  assign wire314 = $signed(wire304[(4'h9):(3'h4)]);
  assign wire315 = $unsigned((~&{$unsigned($signed(wire303)),
                       (^reg311[(1'h0):(1'h0)])}));
  assign wire316 = wire308;
  assign wire317 = {($unsigned($unsigned((8'ha0))) ?
                           (wire310 >> {$unsigned(wire307)}) : wire306)};
  assign wire318 = ($signed(($unsigned(wire315[(5'h10):(2'h3)]) ?
                       ($unsigned((8'hac)) != $unsigned(reg312)) : $signed((|wire306)))) <<< $unsigned((($signed(wire317) <<< (~wire310)) & $unsigned(wire310))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module273
#( parameter param295 = ((!(8'hb5)) ? (~(&(((7'h43) ? (8'hb1) : (8'hbf)) ? ((8'ha1) <= (8'h9f)) : ((7'h43) <= (8'hba))))) : (!(7'h44))) )
(y, clk, wire277, wire276, wire275, wire274);
  output wire [(32'ha7):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire277;
  input wire signed [(5'h10):(1'h0)] wire276;
  input wire signed [(4'ha):(1'h0)] wire275;
  input wire signed [(3'h4):(1'h0)] wire274;
  wire signed [(2'h3):(1'h0)] wire294;
  wire [(4'hf):(1'h0)] wire293;
  wire [(3'h6):(1'h0)] wire292;
  wire [(3'h4):(1'h0)] wire291;
  wire signed [(2'h3):(1'h0)] wire290;
  wire signed [(4'hb):(1'h0)] wire289;
  wire [(4'h9):(1'h0)] wire288;
  wire [(5'h11):(1'h0)] wire287;
  reg [(3'h6):(1'h0)] reg286 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg285 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg284 = (1'h0);
  reg [(5'h11):(1'h0)] reg283 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg282 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg281 = (1'h0);
  reg [(5'h13):(1'h0)] reg280 = (1'h0);
  reg [(2'h2):(1'h0)] reg279 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg278 = (1'h0);
  assign y = {wire294,
                 wire293,
                 wire292,
                 wire291,
                 wire290,
                 wire289,
                 wire288,
                 wire287,
                 reg286,
                 reg285,
                 reg284,
                 reg283,
                 reg282,
                 reg281,
                 reg280,
                 reg279,
                 reg278,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg278 <= {wire277[(4'h8):(3'h6)]};
      if (wire275)
        begin
          reg279 <= (($unsigned(wire277[(4'ha):(1'h0)]) ^~ $signed(((|wire277) ?
                  {wire276, (8'ha7)} : (wire277 || (8'hbe))))) ?
              {($signed(reg278) | wire276),
                  $signed($unsigned((wire274 >>> wire275)))} : wire277);
          if (($unsigned(((((8'hb2) ?
                  reg279 : wire275) == $unsigned(reg279)) || wire275)) ?
              {$signed(((^(8'hb8)) ?
                      (wire275 ?
                          reg279 : wire276) : (!(8'hbe))))} : ((^$signed($signed(wire274))) ?
                  wire277[(1'h0):(1'h0)] : (wire277[(3'h7):(1'h0)] >> ((~|wire274) != (~|(7'h44)))))))
            begin
              reg280 <= wire274[(1'h1):(1'h1)];
              reg281 <= (|reg278[(3'h4):(2'h3)]);
              reg282 <= reg280;
              reg283 <= (({($unsigned((7'h42)) ^~ reg278)} << $signed($unsigned((|wire276)))) ?
                  (~{(~^reg279[(2'h2):(1'h0)])}) : $signed(wire276));
            end
          else
            begin
              reg280 <= (wire276 ?
                  $unsigned(((+(|reg283)) & $signed(((7'h44) ?
                      wire276 : (8'hb0))))) : reg280);
              reg281 <= (~((8'hb1) <<< {reg280}));
              reg282 <= ($unsigned($signed($signed((reg280 ?
                  wire277 : wire277)))) - ($signed($signed($unsigned(wire277))) != {(8'ha1)}));
              reg283 <= ((reg278[(4'hf):(2'h2)] ?
                      wire274 : $unsigned(($unsigned(reg278) != (wire275 >= wire276)))) ?
                  $unsigned($unsigned($unsigned({(8'ha1),
                      (8'hbf)}))) : (^($unsigned((+reg279)) >>> ((8'haa) - wire274[(1'h1):(1'h1)]))));
            end
          reg284 <= ((reg279 ?
              $unsigned($unsigned($unsigned(reg279))) : $signed(($unsigned((8'haf)) ^ reg282))) ~^ (^~{{(~|wire275)},
              ((~|reg280) ? (^~reg278) : reg282[(1'h1):(1'h1)])}));
          reg285 <= (~&(&wire276[(3'h5):(2'h2)]));
          reg286 <= {(reg284 ^~ (~|wire277[(2'h3):(1'h1)]))};
        end
      else
        begin
          reg279 <= $unsigned($unsigned({reg283,
              ((~&reg283) ? $signed((8'hab)) : reg280[(4'hf):(4'hb)])}));
          reg280 <= (!$signed(wire276[(3'h7):(2'h3)]));
          reg281 <= $signed(({reg283[(3'h6):(1'h1)]} ^ ((reg285 & (reg282 ?
              (8'ha0) : wire277)) <= reg280[(4'ha):(2'h3)])));
        end
    end
  assign wire287 = ({(reg283[(4'h9):(3'h7)] == ((&(7'h42)) ?
                               reg280 : (^reg282))),
                           {($unsigned(wire274) ?
                                   (&reg279) : (wire277 ? reg278 : reg279)),
                               (wire276 <<< (8'hae))}} ?
                       reg283 : $signed(((wire276[(3'h6):(3'h5)] ?
                           $signed((8'ha4)) : (~^wire275)) && (((8'hbb) ?
                               reg278 : reg286) ?
                           (reg285 ? wire274 : reg285) : (|wire276)))));
  assign wire288 = ({$signed(((reg282 & wire277) ?
                               (~&reg286) : $unsigned(reg279)))} ?
                       reg282 : $signed(wire277[(4'ha):(3'h5)]));
  assign wire289 = (((reg280 ? $signed($unsigned(reg278)) : {(!(7'h43))}) ?
                           $signed(({reg279} ~^ {wire277,
                               reg281})) : reg282[(4'hb):(4'ha)]) ?
                       (($unsigned((reg282 || wire288)) >> $unsigned($signed(wire274))) ?
                           $signed((-(reg283 ?
                               reg281 : wire274))) : ({$signed(wire274)} ?
                               ({wire287,
                                   wire287} != wire275) : (+$signed(wire275)))) : wire275[(3'h7):(2'h2)]);
  assign wire290 = wire289;
  assign wire291 = reg282[(3'h7):(1'h1)];
  assign wire292 = (~|reg285[(1'h0):(1'h0)]);
  assign wire293 = {({$signed($unsigned(wire276))} ?
                           ($unsigned({reg282}) ?
                               $signed($unsigned(wire277)) : ($signed(reg282) ?
                                   reg279 : (reg278 ?
                                       reg284 : wire292))) : wire292)};
  assign wire294 = $unsigned($signed((|($unsigned(wire293) * reg284[(1'h1):(1'h0)]))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module252
#(parameter param266 = (8'haa), parameter param267 = param266)
(y, clk, wire256, wire255, wire254, wire253);
  output wire [(32'h75):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire256;
  input wire signed [(4'hf):(1'h0)] wire255;
  input wire signed [(4'hd):(1'h0)] wire254;
  input wire [(5'h11):(1'h0)] wire253;
  wire signed [(2'h2):(1'h0)] wire265;
  wire [(4'he):(1'h0)] wire264;
  wire [(5'h15):(1'h0)] wire263;
  wire [(3'h5):(1'h0)] wire262;
  wire signed [(5'h10):(1'h0)] wire261;
  wire signed [(4'hd):(1'h0)] wire260;
  wire [(3'h5):(1'h0)] wire259;
  wire [(5'h14):(1'h0)] wire258;
  wire [(5'h14):(1'h0)] wire257;
  assign y = {wire265,
                 wire264,
                 wire263,
                 wire262,
                 wire261,
                 wire260,
                 wire259,
                 wire258,
                 wire257,
                 (1'h0)};
  assign wire257 = (wire254 & wire253);
  assign wire258 = $unsigned($signed(wire254[(3'h6):(2'h3)]));
  assign wire259 = wire258;
  assign wire260 = (|wire259[(3'h4):(1'h1)]);
  assign wire261 = (((wire253 && {{wire256, wire258}, $signed(wire260)}) ?
                       wire258[(3'h4):(2'h2)] : wire257) != ($signed(wire255[(4'hc):(2'h2)]) ?
                       (8'hae) : wire258[(4'h9):(3'h5)]));
  assign wire262 = ($unsigned($signed($unsigned((wire257 ?
                           wire259 : wire257)))) ?
                       $signed((8'ha8)) : {wire253});
  assign wire263 = wire257;
  assign wire264 = wire259[(1'h1):(1'h1)];
  assign wire265 = ($unsigned(($signed($signed(wire259)) ?
                           $unsigned($signed(wire257)) : wire258)) ?
                       (^~$signed($signed((wire259 || wire262)))) : $unsigned({{wire259,
                               {wire258, wire254}},
                           wire260[(4'h9):(3'h4)]}));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module203
#( parameter param224 = (({(-((8'h9f) ? (8'h9d) : (8'ha9))), (((7'h41) && (8'hb9)) ? (^~(8'hb4)) : {(7'h40), (8'hb5)})} ? ({((8'haa) <<< (8'ha7))} >= ({(8'haf)} ? ((8'ha8) ? (8'ha5) : (8'h9e)) : (^(8'ha1)))) : (^((&(8'hb8)) - ((8'ha8) ? (8'hbb) : (8'hae))))) ? (^~(((+(8'hac)) ? ((8'hb4) && (8'h9e)) : ((8'hb4) ? (8'haf) : (8'ha5))) ? ((!(8'hba)) ? ((8'ha1) ? (8'hae) : (8'hbe)) : {(8'hb0), (8'hb9)}) : {((8'hab) ? (8'h9c) : (8'hbc)), ((8'ha0) ? (8'hb5) : (8'hb3))})) : (-{(((8'haf) ? (8'hb5) : (8'ha5)) ~^ (~&(8'ha8)))}))
, parameter param225 = ((-(~|param224)) > param224) )
(y, clk, wire208, wire207, wire206, wire205, wire204);
  output wire [(32'h95):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h7):(1'h0)] wire208;
  input wire signed [(4'ha):(1'h0)] wire207;
  input wire [(3'h5):(1'h0)] wire206;
  input wire signed [(5'h11):(1'h0)] wire205;
  input wire signed [(4'he):(1'h0)] wire204;
  wire signed [(2'h3):(1'h0)] wire223;
  wire [(4'hb):(1'h0)] wire222;
  wire [(4'h8):(1'h0)] wire221;
  wire signed [(3'h6):(1'h0)] wire220;
  wire signed [(3'h7):(1'h0)] wire219;
  wire signed [(5'h15):(1'h0)] wire218;
  wire signed [(4'h8):(1'h0)] wire217;
  wire [(4'ha):(1'h0)] wire216;
  wire [(4'hb):(1'h0)] wire215;
  wire signed [(2'h2):(1'h0)] wire214;
  wire [(3'h7):(1'h0)] wire213;
  wire [(4'hd):(1'h0)] wire212;
  wire [(5'h12):(1'h0)] wire211;
  wire [(2'h2):(1'h0)] wire210;
  wire signed [(5'h15):(1'h0)] wire209;
  assign y = {wire223,
                 wire222,
                 wire221,
                 wire220,
                 wire219,
                 wire218,
                 wire217,
                 wire216,
                 wire215,
                 wire214,
                 wire213,
                 wire212,
                 wire211,
                 wire210,
                 wire209,
                 (1'h0)};
  assign wire209 = ($signed($signed($unsigned(((8'h9f) ? wire204 : (7'h41))))) ?
                       (((~^(wire206 ? wire204 : wire205)) ?
                           (~&wire207[(2'h2):(1'h1)]) : (~&$signed(wire204))) > {$signed((wire205 ?
                               wire205 : wire207)),
                           $signed((wire207 ^ wire204))}) : (~^($signed(wire204[(4'ha):(4'h8)]) ~^ wire206)));
  assign wire210 = ($unsigned((8'hb5)) ?
                       $signed($unsigned({(wire208 ^ wire208)})) : ((-wire205) ?
                           {((wire209 || (8'ha4)) < wire209),
                               $signed($unsigned(wire206))} : $signed((&(wire204 ~^ wire209)))));
  assign wire211 = $unsigned($unsigned(((^(~|wire208)) >= wire204[(2'h3):(1'h0)])));
  assign wire212 = $unsigned(wire208[(2'h3):(2'h2)]);
  assign wire213 = wire208[(3'h6):(3'h4)];
  assign wire214 = (wire207[(4'ha):(4'ha)] ? wire209 : (8'hb6));
  assign wire215 = wire207;
  assign wire216 = $signed((wire212[(4'hc):(2'h3)] ?
                       {((wire208 ? wire211 : wire213) ?
                               $unsigned(wire205) : (wire212 == wire209)),
                           $unsigned($signed(wire210))} : (~({(8'ha2),
                               wire204} ?
                           wire210 : (wire207 ? wire215 : (8'hb3))))));
  assign wire217 = (~($signed(wire205) ^ $unsigned($unsigned($signed(wire216)))));
  assign wire218 = wire211;
  assign wire219 = {(wire207 ?
                           ($signed($unsigned((8'had))) ?
                               {wire204[(4'hd):(3'h4)],
                                   (wire211 * wire205)} : {(wire206 <<< wire217)}) : wire212[(3'h7):(3'h7)]),
                       $signed($unsigned((|(wire211 != wire214))))};
  assign wire220 = ($signed(wire210) ?
                       $signed((-(~|$signed(wire208)))) : ($signed((-(wire219 >>> (8'hb3)))) < wire217[(3'h4):(2'h3)]));
  assign wire221 = (!($unsigned(wire208) + wire210[(1'h1):(1'h1)]));
  assign wire222 = $signed(wire210);
  assign wire223 = ({wire220, (wire218 >>> wire222)} & $unsigned(wire210));
endmodule