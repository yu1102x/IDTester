(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param185 = (~(8'haa)))
(y, clk, wire0, wire1, wire2, wire3);
  output wire [(32'hbe):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h2):(1'h0)] wire0;
  input wire signed [(5'h13):(1'h0)] wire1;
  input wire signed [(5'h14):(1'h0)] wire2;
  input wire [(5'h15):(1'h0)] wire3;
  wire signed [(4'h9):(1'h0)] wire184;
  wire signed [(3'h4):(1'h0)] wire183;
  wire signed [(5'h14):(1'h0)] wire182;
  wire signed [(4'ha):(1'h0)] wire181;
  wire signed [(5'h11):(1'h0)] wire4;
  wire signed [(5'h14):(1'h0)] wire5;
  wire [(4'hc):(1'h0)] wire6;
  wire [(5'h12):(1'h0)] wire170;
  wire [(3'h7):(1'h0)] wire172;
  reg signed [(4'h8):(1'h0)] reg173 = (1'h0);
  reg [(4'ha):(1'h0)] reg174 = (1'h0);
  wire [(3'h4):(1'h0)] wire175;
  reg signed [(4'h9):(1'h0)] reg176 = (1'h0);
  wire [(3'h7):(1'h0)] wire177;
  wire signed [(5'h14):(1'h0)] wire178;
  wire signed [(4'he):(1'h0)] wire179;
  assign y = {wire184,
                 wire183,
                 wire182,
                 wire181,
                 wire4,
                 wire5,
                 wire6,
                 wire170,
                 wire172,
                 reg173,
                 reg174,
                 wire175,
                 reg176,
                 wire177,
                 wire178,
                 wire179,
                 (1'h0)};
  assign wire4 = wire2;
  assign wire5 = wire3[(2'h2):(2'h2)];
  assign wire6 = wire2;
  module7 modinst171 (.wire11(wire6), .wire10(wire2), .wire9(wire1), .clk(clk), .wire8(wire5), .y(wire170));
  assign wire172 = (($unsigned(wire0[(2'h2):(1'h1)]) ^ (wire3[(5'h14):(5'h14)] ?
                       (!(wire6 <<< wire170)) : wire170)) * (&$signed(wire3[(5'h10):(4'ha)])));
  always
    @(posedge clk) begin
      reg173 <= $signed($unsigned(((&(wire5 <<< wire4)) >= (~$unsigned((8'hb9))))));
    end
  always
    @(posedge clk) begin
      reg174 <= wire2[(3'h4):(3'h4)];
    end
  assign wire175 = wire1;
  always
    @(posedge clk) begin
      reg176 <= ((|{$unsigned((wire0 & wire2)),
          wire1[(5'h10):(3'h4)]}) != (^~$signed($signed($unsigned(wire172)))));
    end
  assign wire177 = $unsigned($signed((~|(8'ha0))));
  assign wire178 = wire177;
  module56 modinst180 (.y(wire179), .clk(clk), .wire61(wire3), .wire58(reg174), .wire60(wire4), .wire57(reg176), .wire59(wire178));
  assign wire181 = $unsigned($signed(wire170));
  assign wire182 = (((wire3[(4'hd):(1'h0)] ?
                           {$signed(wire0), (wire1 > reg176)} : (-(^(8'hac)))) ?
                       $unsigned($signed(wire6[(4'h9):(1'h1)])) : (((&wire4) ~^ wire170) ?
                           (!(~|wire4)) : wire170[(4'h9):(4'h8)])) && ($unsigned(reg173) >> (~&((wire175 - wire179) >>> {(8'hbf)}))));
  assign wire183 = $signed({$signed(((wire1 + reg173) ?
                           wire3[(2'h3):(2'h3)] : reg176[(1'h1):(1'h0)])),
                       wire170[(1'h0):(1'h0)]});
  assign wire184 = (~wire181);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module7
#( parameter param169 = {((((~|(8'ha2)) ? ((8'hbc) < (8'ha2)) : ((8'ha8) ? (8'haf) : (7'h44))) ? (|(8'h9d)) : {(8'h9e), {(8'hb6), (8'hb5)}}) ^~ {(~|((8'ha6) ? (8'hbe) : (8'ha7)))})} )
(y, clk, wire8, wire9, wire10, wire11);
  output wire [(32'h189):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire8;
  input wire [(5'h13):(1'h0)] wire9;
  input wire signed [(5'h13):(1'h0)] wire10;
  input wire [(4'hc):(1'h0)] wire11;
  wire signed [(5'h13):(1'h0)] wire168;
  reg signed [(5'h15):(1'h0)] reg167 = (1'h0);
  reg [(4'h9):(1'h0)] reg166 = (1'h0);
  reg [(5'h14):(1'h0)] reg165 = (1'h0);
  reg signed [(4'he):(1'h0)] reg164 = (1'h0);
  reg signed [(4'he):(1'h0)] reg163 = (1'h0);
  reg [(4'hd):(1'h0)] reg162 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg161 = (1'h0);
  reg [(5'h10):(1'h0)] reg160 = (1'h0);
  wire [(3'h7):(1'h0)] wire159;
  wire signed [(3'h6):(1'h0)] wire158;
  wire [(5'h13):(1'h0)] wire156;
  wire [(4'hb):(1'h0)] wire155;
  wire [(4'he):(1'h0)] wire154;
  reg [(4'h8):(1'h0)] reg153 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire152;
  wire signed [(3'h6):(1'h0)] wire151;
  wire [(3'h7):(1'h0)] wire82;
  wire signed [(5'h15):(1'h0)] wire55;
  wire [(4'hd):(1'h0)] wire54;
  wire signed [(4'hb):(1'h0)] wire12;
  wire signed [(4'ha):(1'h0)] wire30;
  wire signed [(5'h14):(1'h0)] wire52;
  wire signed [(5'h11):(1'h0)] wire84;
  wire signed [(5'h14):(1'h0)] wire85;
  wire [(5'h13):(1'h0)] wire86;
  wire signed [(5'h12):(1'h0)] wire87;
  wire [(4'hb):(1'h0)] wire136;
  wire [(3'h7):(1'h0)] wire149;
  assign y = {wire168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 wire159,
                 wire158,
                 wire156,
                 wire155,
                 wire154,
                 reg153,
                 wire152,
                 wire151,
                 wire82,
                 wire55,
                 wire54,
                 wire12,
                 wire30,
                 wire52,
                 wire84,
                 wire85,
                 wire86,
                 wire87,
                 wire136,
                 wire149,
                 (1'h0)};
  assign wire12 = wire10;
  module13 modinst31 (wire30, clk, wire8, wire9, wire12, wire10);
  module32 modinst53 (wire52, clk, wire9, wire11, wire10, wire30, wire12);
  assign wire54 = wire9;
  assign wire55 = $signed(((|(8'ha2)) ?
                      $unsigned($signed($signed(wire9))) : (wire54[(4'h8):(4'h8)] ?
                          wire8 : $unsigned({wire54}))));
  module56 modinst83 (wire82, clk, wire10, wire55, wire52, wire30, wire8);
  assign wire84 = wire9;
  assign wire85 = {wire82,
                      (((8'h9e) - (wire12 - wire52)) ?
                          (~^(wire8 ?
                              $unsigned(wire55) : (^~wire84))) : $signed($unsigned(wire11)))};
  assign wire86 = $signed((+((!(wire8 ^~ (8'haf))) & wire55)));
  assign wire87 = $unsigned($signed($signed(wire82[(3'h6):(3'h6)])));
  module88 modinst137 (.wire90(wire11), .y(wire136), .wire89(wire8), .clk(clk), .wire91(wire84), .wire92(wire52));
  module138 modinst150 (.wire140(wire55), .y(wire149), .wire139(wire84), .wire141(wire54), .wire143(wire9), .clk(clk), .wire142(wire85));
  assign wire151 = wire10[(4'he):(3'h4)];
  assign wire152 = (!wire87[(4'hf):(1'h0)]);
  always
    @(posedge clk) begin
      reg153 <= $unsigned((^$signed(((~|wire85) ?
          ((8'ha2) <<< wire149) : $signed(wire8)))));
    end
  assign wire154 = wire8;
  assign wire155 = ($signed(($signed((wire10 & (8'hb2))) ?
                       wire84[(4'ha):(4'h8)] : ((~(7'h43)) ?
                           $unsigned(wire84) : (wire87 != wire10)))) ^~ wire154[(3'h6):(2'h2)]);
  module88 modinst157 (wire156, clk, wire155, wire136, wire86, wire54);
  assign wire158 = (~&((({wire154} ? (wire82 ? wire52 : wire82) : (&(8'ha6))) ?
                           {(wire86 < wire156)} : {(wire10 <= wire85),
                               wire12[(3'h7):(1'h0)]}) ?
                       wire11[(4'ha):(2'h2)] : $signed($unsigned(wire8))));
  assign wire159 = {({wire151[(1'h0):(1'h0)]} <= (wire55[(5'h11):(3'h6)] ^~ $signed(((7'h43) ?
                           wire87 : wire10)))),
                       $signed($unsigned(($unsigned(wire10) + $unsigned(wire86))))};
  always
    @(posedge clk) begin
      reg160 <= wire158[(3'h4):(2'h3)];
      if ({({(-wire52)} ?
              $signed(((wire158 ?
                  wire11 : wire55) & wire9[(5'h10):(3'h4)])) : $unsigned(wire151)),
          ($signed((wire9[(4'hf):(3'h5)] >> ((8'ha2) ? wire156 : wire85))) ?
              ({$signed(wire156), ((8'hb5) ? wire9 : wire87)} ?
                  ({(8'ha5)} ?
                      (|wire30) : (~&wire54)) : (wire86[(5'h11):(4'hb)] == wire84)) : wire82[(1'h0):(1'h0)])})
        begin
          reg161 <= wire12;
          reg162 <= $unsigned(wire84);
          reg163 <= wire84[(4'hc):(1'h1)];
          if (reg153[(1'h0):(1'h0)])
            begin
              reg164 <= (&(8'ha4));
              reg165 <= $unsigned({$signed(($unsigned(wire152) + wire11[(4'h9):(3'h5)]))});
            end
          else
            begin
              reg164 <= ((($unsigned($unsigned(wire156)) & wire158[(2'h2):(1'h1)]) ^ $signed(reg164)) ?
                  (reg153 ?
                      (^~(~(reg162 ?
                          wire84 : reg165))) : ({reg163[(3'h4):(1'h0)]} ?
                          wire86[(5'h12):(4'hd)] : ((!reg160) & (wire87 < reg161)))) : (reg160 << wire82[(1'h1):(1'h0)]));
              reg165 <= {reg161};
              reg166 <= $unsigned(wire84[(2'h3):(1'h1)]);
              reg167 <= wire151[(1'h1):(1'h0)];
            end
        end
      else
        begin
          reg161 <= $unsigned($signed((^(-wire11[(1'h0):(1'h0)]))));
          reg162 <= (wire84 ?
              ((~^{(wire136 ? wire87 : reg165)}) ?
                  wire82[(2'h3):(2'h3)] : $signed(($signed(wire155) ?
                      wire151 : ((8'ha1) ~^ wire54)))) : (wire156 | wire86[(4'h8):(3'h6)]));
          if ((|(({(wire87 | wire155)} ^~ (+(wire155 ? wire54 : wire9))) ?
              $unsigned(((~^wire11) ?
                  $signed(wire12) : (^~reg166))) : (~|((wire154 ?
                      wire156 : reg163) ?
                  $unsigned(wire87) : (~|wire82))))))
            begin
              reg163 <= $signed($unsigned((^~(-{wire11}))));
              reg164 <= $unsigned(wire87[(3'h4):(1'h0)]);
              reg165 <= $unsigned(wire85[(4'ha):(1'h0)]);
            end
          else
            begin
              reg163 <= (^~{({reg160[(4'ha):(2'h3)]} ^ $unsigned((wire12 | wire151)))});
              reg164 <= (^~wire156);
              reg165 <= wire11;
              reg166 <= reg163;
              reg167 <= (+(wire30 ?
                  $unsigned({$unsigned((7'h41))}) : {wire54[(3'h4):(2'h3)]}));
            end
        end
    end
  assign wire168 = (|((~|(~&{wire11,
                       wire11})) - (($unsigned(wire158) > ((8'haa) ?
                           reg166 : reg161)) ?
                       reg160[(4'he):(1'h1)] : (+wire12))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module138  (y, clk, wire143, wire142, wire141, wire140, wire139);
  output wire [(32'h34):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'he):(1'h0)] wire143;
  input wire [(5'h11):(1'h0)] wire142;
  input wire signed [(4'h8):(1'h0)] wire141;
  input wire signed [(5'h15):(1'h0)] wire140;
  input wire signed [(5'h10):(1'h0)] wire139;
  wire [(4'ha):(1'h0)] wire148;
  wire signed [(3'h7):(1'h0)] wire147;
  wire [(3'h5):(1'h0)] wire146;
  wire signed [(4'hb):(1'h0)] wire145;
  wire [(5'h12):(1'h0)] wire144;
  assign y = {wire148, wire147, wire146, wire145, wire144, (1'h0)};
  assign wire144 = $signed(((wire140 ?
                       {$unsigned((7'h44)),
                           (wire142 ?
                               wire143 : wire141)} : wire142[(3'h6):(3'h5)]) <= $signed(wire141)));
  assign wire145 = (8'ha8);
  assign wire146 = $unsigned((((7'h43) ?
                           $unsigned((wire141 <= wire144)) : ($unsigned(wire142) ?
                               $unsigned(wire140) : wire140)) ?
                       wire139[(4'he):(1'h0)] : wire145[(4'hb):(3'h4)]));
  assign wire147 = wire146[(1'h1):(1'h1)];
  assign wire148 = ((wire140 >= ($signed(((8'hb9) ? wire147 : wire140)) ?
                       ($signed(wire147) ?
                           (wire146 ?
                               wire142 : wire145) : (wire142 == wire139)) : (wire141[(1'h1):(1'h1)] - wire140))) == wire143[(1'h0):(1'h0)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module88
#( parameter param135 = ((|(((^(8'h9f)) ? (|(8'ha9)) : (8'hb6)) << (~|(~^(8'hb7))))) ? ((!(!(+(8'hb9)))) ? (-(~^((8'hb3) && (8'hbd)))) : ({{(8'ha6)}} != (~&((8'ha7) ? (8'hb7) : (8'hbf))))) : ((8'ha8) ? ((((8'hb3) < (8'ha5)) == ((8'ha7) ? (8'hb2) : (8'hbd))) ? (^((8'ha2) ? (8'hb9) : (8'haa))) : {{(8'ha9), (8'ha5)}, (+(8'h9e))}) : ({(~^(8'h9f))} >> ((~^(8'hab)) >> ((7'h44) <= (8'hb1)))))) )
(y, clk, wire92, wire91, wire90, wire89);
  output wire [(32'h1f9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire92;
  input wire signed [(2'h2):(1'h0)] wire91;
  input wire signed [(4'ha):(1'h0)] wire90;
  input wire signed [(4'h8):(1'h0)] wire89;
  reg [(2'h3):(1'h0)] reg134 = (1'h0);
  reg [(5'h15):(1'h0)] reg133 = (1'h0);
  reg [(3'h4):(1'h0)] reg132 = (1'h0);
  reg [(4'he):(1'h0)] reg131 = (1'h0);
  reg [(4'hd):(1'h0)] reg130 = (1'h0);
  reg [(4'h8):(1'h0)] reg129 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg128 = (1'h0);
  reg [(4'ha):(1'h0)] reg127 = (1'h0);
  reg [(3'h4):(1'h0)] reg126 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg125 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg124 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg123 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg122 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg121 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg120 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg119 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire118;
  wire [(4'h8):(1'h0)] wire117;
  reg signed [(5'h14):(1'h0)] reg116 = (1'h0);
  reg [(5'h14):(1'h0)] reg115 = (1'h0);
  reg [(4'hb):(1'h0)] reg114 = (1'h0);
  reg [(4'ha):(1'h0)] reg113 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire112;
  wire signed [(4'ha):(1'h0)] wire111;
  wire signed [(5'h11):(1'h0)] wire110;
  wire [(5'h10):(1'h0)] wire109;
  wire signed [(5'h12):(1'h0)] wire108;
  wire [(4'ha):(1'h0)] wire107;
  wire [(5'h10):(1'h0)] wire106;
  wire signed [(4'h8):(1'h0)] wire105;
  wire [(5'h12):(1'h0)] wire104;
  wire [(5'h15):(1'h0)] wire103;
  wire signed [(5'h11):(1'h0)] wire102;
  wire signed [(4'h8):(1'h0)] wire101;
  wire signed [(4'ha):(1'h0)] wire100;
  reg signed [(4'h8):(1'h0)] reg99 = (1'h0);
  reg [(4'ha):(1'h0)] reg98 = (1'h0);
  reg [(3'h6):(1'h0)] reg97 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg96 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg95 = (1'h0);
  reg [(5'h13):(1'h0)] reg94 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg93 = (1'h0);
  assign y = {reg134,
                 reg133,
                 reg132,
                 reg131,
                 reg130,
                 reg129,
                 reg128,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 reg121,
                 reg120,
                 reg119,
                 wire118,
                 wire117,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 wire112,
                 wire111,
                 wire110,
                 wire109,
                 wire108,
                 wire107,
                 wire106,
                 wire105,
                 wire104,
                 wire103,
                 wire102,
                 wire101,
                 wire100,
                 reg99,
                 reg98,
                 reg97,
                 reg96,
                 reg95,
                 reg94,
                 reg93,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg93 <= wire89[(4'h8):(4'h8)];
      if (wire90[(1'h0):(1'h0)])
        begin
          reg94 <= (!($unsigned(({wire89, wire91} ?
              $unsigned(wire90) : (&wire92))) << $signed(($unsigned(wire91) <= ((8'ha2) ?
              (7'h42) : wire92)))));
          reg95 <= (^($signed($signed($signed(reg94))) ?
              (+$signed((wire90 ? wire91 : reg93))) : wire91));
          reg96 <= wire89[(3'h5):(3'h5)];
          reg97 <= $signed((|wire91[(2'h2):(2'h2)]));
        end
      else
        begin
          reg94 <= (~$signed(wire91[(1'h0):(1'h0)]));
          if (((wire92 ~^ $signed(($unsigned(reg96) ?
              reg97 : $unsigned(wire89)))) != wire92))
            begin
              reg95 <= ((wire91 != ((-reg95[(3'h7):(2'h2)]) ~^ (^~((8'hb1) ?
                  reg93 : (8'hbc))))) ~^ ($signed(reg97[(1'h0):(1'h0)]) ?
                  (((reg95 ?
                      (8'hab) : reg94) >= $signed(reg95)) << wire90[(2'h2):(2'h2)]) : ($signed((8'hb1)) ?
                      reg95[(3'h4):(1'h1)] : $signed((^wire91)))));
            end
          else
            begin
              reg95 <= (&$unsigned(reg93));
              reg96 <= wire89[(3'h4):(2'h2)];
              reg97 <= (!reg96);
            end
          reg98 <= (^$unsigned(wire90));
        end
      reg99 <= (|{reg96[(1'h0):(1'h0)], (reg98 ? wire92 : wire92)});
    end
  assign wire100 = {$signed($unsigned(reg99[(1'h1):(1'h1)])),
                       $signed(((((8'hb1) <= reg99) <= (wire91 ?
                           reg97 : reg94)) >= $unsigned((+(8'ha7)))))};
  assign wire101 = reg99;
  assign wire102 = $unsigned((^reg96));
  assign wire103 = wire100;
  assign wire104 = $unsigned((~^((8'hba) & reg95)));
  assign wire105 = $signed(({wire89[(3'h5):(2'h2)],
                       reg97} ^~ {$unsigned(wire102[(2'h2):(2'h2)]),
                       $unsigned($unsigned(reg97))}));
  assign wire106 = ((7'h41) ?
                       wire89[(2'h3):(2'h2)] : (reg97[(3'h4):(1'h1)] ?
                           (reg99 ?
                               {wire100} : {{reg97, reg93}, (8'hb3)}) : reg99));
  assign wire107 = $unsigned((~&$unsigned({(reg97 ? (8'hbf) : reg97)})));
  assign wire108 = (+reg97[(3'h6):(3'h6)]);
  assign wire109 = reg98;
  assign wire110 = (~(wire107 ?
                       ({(wire89 ? reg98 : reg98),
                           {wire105,
                               wire89}} < (+(~^(7'h40)))) : {reg99[(2'h3):(1'h1)],
                           ($signed(wire90) < $unsigned(reg97))}));
  assign wire111 = (|$signed(($signed($signed(reg94)) ^ $unsigned($unsigned(wire110)))));
  assign wire112 = (($unsigned(wire102[(3'h4):(2'h2)]) ?
                       wire105[(4'h8):(3'h4)] : (wire110 ?
                           $unsigned($unsigned(reg93)) : ((-(8'ha8)) ?
                               wire102[(1'h0):(1'h0)] : wire102[(1'h1):(1'h0)]))) >>> wire111);
  always
    @(posedge clk) begin
      reg113 <= $unsigned($unsigned($signed(($unsigned((8'hb3)) ?
          wire90[(3'h4):(2'h2)] : (~^(8'hb7))))));
      reg114 <= $unsigned({((~$unsigned(reg97)) ?
              $unsigned((wire100 ? wire103 : (8'hb3))) : ($signed(wire89) ?
                  wire109 : (8'hab))),
          wire106[(3'h7):(2'h3)]});
      reg115 <= reg96[(2'h2):(1'h0)];
      reg116 <= $unsigned((~wire108[(5'h10):(2'h3)]));
    end
  assign wire117 = $unsigned({(($signed(wire107) ?
                           wire112 : (wire101 ?
                               wire103 : wire105)) >>> ($signed((8'h9f)) ?
                           (reg93 < reg97) : (8'haf))),
                       wire111[(3'h4):(2'h3)]});
  assign wire118 = (8'hb7);
  always
    @(posedge clk) begin
      if ((($signed($unsigned((wire91 ?
          wire104 : wire103))) >= $signed(((wire92 <= wire100) || (8'hb6)))) >= wire103))
        begin
          reg119 <= (($unsigned({wire100[(2'h2):(1'h1)],
                  {wire109}}) ~^ ($unsigned((reg94 ^ wire106)) ?
                  reg98 : ((~&(8'hbd)) ?
                      reg93[(3'h4):(1'h1)] : $unsigned(wire105)))) ?
              $unsigned($unsigned(({reg114} | $unsigned(reg116)))) : (8'ha6));
          if ($unsigned((((~(wire117 & wire103)) ?
                  (reg113[(1'h1):(1'h0)] ?
                      $signed((8'ha3)) : {(7'h44)}) : $signed($unsigned(wire111))) ?
              $signed((8'hbc)) : ($signed($signed(wire111)) ?
                  wire90 : wire107))))
            begin
              reg120 <= reg95[(4'ha):(3'h7)];
              reg121 <= (((~$signed($signed(wire100))) ?
                  (($unsigned(wire89) > (reg97 ? wire109 : wire108)) ?
                      $unsigned(wire104[(5'h11):(3'h5)]) : ((~&reg120) ~^ wire117)) : $unsigned((reg113[(3'h4):(1'h0)] ?
                      {reg97,
                          (8'hbb)} : (^(8'ha8))))) - (^~$unsigned($unsigned($unsigned(wire102)))));
              reg122 <= (wire117[(3'h4):(3'h4)] * reg96);
            end
          else
            begin
              reg120 <= $unsigned(((&(~^(wire100 << reg115))) & (($unsigned(wire112) || $unsigned(wire104)) ?
                  wire100[(3'h5):(1'h0)] : wire109[(3'h4):(2'h3)])));
            end
          reg123 <= ({($unsigned(((8'h9c) ? reg120 : reg98)) <= reg113)} ?
              $signed(wire100[(4'h9):(3'h7)]) : reg115[(4'hc):(3'h4)]);
          reg124 <= $signed(reg123);
        end
      else
        begin
          reg119 <= ($signed({(!wire106[(2'h3):(1'h0)])}) >>> (^$signed($unsigned(reg94))));
          reg120 <= $unsigned({(8'hae)});
          reg121 <= (~(~($signed({reg93}) ?
              (reg99 ?
                  $unsigned(reg116) : (reg116 << wire111)) : (-{wire111}))));
          if (wire111)
            begin
              reg122 <= ($unsigned(reg124) <<< (~|((8'ha9) || {(wire106 ?
                      reg98 : wire100)})));
              reg123 <= $unsigned(reg124);
            end
          else
            begin
              reg122 <= ($signed(reg94[(4'hf):(4'h9)]) ?
                  $unsigned(wire106) : (|($signed(wire91) >>> $unsigned($unsigned(reg115)))));
              reg123 <= {wire92[(3'h6):(1'h1)]};
            end
        end
      reg125 <= reg97[(1'h1):(1'h1)];
      if ({(8'hb7)})
        begin
          reg126 <= ($unsigned((($unsigned(reg122) ?
                      {reg95} : wire105[(2'h3):(1'h1)]) ?
                  $unsigned(wire104[(3'h5):(2'h2)]) : $signed(reg98[(3'h4):(1'h0)]))) ?
              $signed((|(+(reg114 ?
                  (8'ha5) : wire89)))) : (reg113[(4'h8):(3'h4)] ?
                  wire101 : (~^$unsigned((~|wire104)))));
          reg127 <= $signed(wire112[(1'h1):(1'h1)]);
          reg128 <= (!reg122[(4'hb):(2'h3)]);
        end
      else
        begin
          reg126 <= (($signed($unsigned((reg116 ?
              wire102 : wire91))) == reg116[(4'h8):(3'h4)]) | (reg114[(4'ha):(3'h6)] ?
              reg126[(1'h0):(1'h0)] : wire90[(3'h4):(2'h2)]));
          if (reg121)
            begin
              reg127 <= (((&(~&$signed(reg95))) ?
                  ({(|wire103), wire91[(1'h0):(1'h0)]} ?
                      ({wire108} - {reg125,
                          wire89}) : (-$unsigned(wire107))) : {$unsigned(((8'hbb) ^ wire109)),
                      {reg121[(1'h1):(1'h1)],
                          (reg94 ?
                              wire103 : reg114)}}) <= (($signed(wire100[(4'h9):(2'h3)]) ?
                  $signed($unsigned(wire107)) : (reg125 ?
                      (~(8'ha8)) : wire117)) ~^ $signed((~|(~(7'h44))))));
              reg128 <= ($unsigned({$signed((reg124 < (8'hb1)))}) ^ $signed(($signed(reg113[(1'h1):(1'h1)]) & (^$signed(wire91)))));
            end
          else
            begin
              reg127 <= wire112[(4'he):(4'hd)];
              reg128 <= $signed($unsigned(reg96[(1'h1):(1'h0)]));
            end
          if (($signed(({wire91[(2'h2):(2'h2)]} ?
                  $unsigned((wire111 > (8'ha7))) : {$unsigned(wire118)})) ?
              {wire101} : $signed(wire110)))
            begin
              reg129 <= $signed((^~(&$unsigned(wire103))));
              reg130 <= $unsigned(wire106);
              reg131 <= $signed($unsigned(((reg113 == $unsigned(wire90)) ?
                  (^reg93) : $signed((!reg114)))));
              reg132 <= reg113;
              reg133 <= (^~(8'hbd));
            end
          else
            begin
              reg129 <= {{reg131}};
              reg130 <= (^~(^(($signed(wire105) ?
                  reg98[(1'h0):(1'h0)] : wire111) - wire108)));
              reg131 <= (~(^(~|reg130)));
            end
        end
      reg134 <= wire100;
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module56
#( parameter param80 = ((^~((((8'hbd) ^ (8'hb2)) != {(8'ha4)}) ? (((8'had) < (8'hb2)) >> (+(8'hbf))) : (~&((8'hb2) | (8'hb2))))) == ((^~(^((8'hb1) < (8'hbb)))) >>> ({(+(8'ha4))} * (8'h9c))))
, parameter param81 = param80 )
(y, clk, wire61, wire60, wire59, wire58, wire57);
  output wire [(32'h97):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire61;
  input wire [(4'he):(1'h0)] wire60;
  input wire [(5'h14):(1'h0)] wire59;
  input wire [(4'ha):(1'h0)] wire58;
  input wire [(4'h9):(1'h0)] wire57;
  wire [(5'h11):(1'h0)] wire79;
  reg signed [(5'h10):(1'h0)] reg78 = (1'h0);
  reg [(2'h2):(1'h0)] reg77 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg76 = (1'h0);
  reg [(4'hf):(1'h0)] reg75 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg74 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg73 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire72;
  wire signed [(2'h2):(1'h0)] wire71;
  wire [(4'ha):(1'h0)] wire70;
  wire signed [(3'h6):(1'h0)] wire69;
  wire signed [(3'h4):(1'h0)] wire68;
  wire signed [(4'h9):(1'h0)] wire67;
  wire signed [(3'h5):(1'h0)] wire66;
  wire signed [(3'h5):(1'h0)] wire65;
  wire signed [(4'h8):(1'h0)] wire64;
  wire [(3'h4):(1'h0)] wire63;
  wire signed [(4'hf):(1'h0)] wire62;
  assign y = {wire79,
                 reg78,
                 reg77,
                 reg76,
                 reg75,
                 reg74,
                 reg73,
                 wire72,
                 wire71,
                 wire70,
                 wire69,
                 wire68,
                 wire67,
                 wire66,
                 wire65,
                 wire64,
                 wire63,
                 wire62,
                 (1'h0)};
  assign wire62 = wire61;
  assign wire63 = $signed((wire57 + $signed($unsigned((wire62 <= wire61)))));
  assign wire64 = ($unsigned(wire57) ^ wire59);
  assign wire65 = $unsigned((-(wire63 ?
                      $signed(wire63[(2'h2):(1'h0)]) : (wire64 * (~wire59)))));
  assign wire66 = wire58;
  assign wire67 = wire58[(1'h0):(1'h0)];
  assign wire68 = (8'ha9);
  assign wire69 = (wire61[(2'h3):(1'h1)] ?
                      (8'hbe) : $signed($signed($signed(wire59))));
  assign wire70 = (wire68 ?
                      ($signed({wire68}) ?
                          ({wire66[(2'h2):(2'h2)]} ?
                              {wire61} : $signed(wire61[(2'h3):(2'h2)])) : $signed($unsigned(wire69[(1'h0):(1'h0)]))) : ((wire64[(2'h2):(2'h2)] ?
                              (^~(wire69 ^~ wire60)) : $unsigned((&wire63))) ?
                          wire61 : wire67));
  assign wire71 = ($signed($signed($signed((^~wire59)))) + $signed($unsigned($signed($unsigned((7'h43))))));
  assign wire72 = ((~^$signed((+wire68))) == (wire69 ^~ ($unsigned((~^(8'h9f))) ?
                      wire71 : $signed((wire63 ? wire59 : wire69)))));
  always
    @(posedge clk) begin
      if ((wire64[(3'h5):(2'h2)] <= ((($unsigned(wire71) >> $signed(wire59)) + $signed($unsigned((7'h44)))) ?
          $signed((wire65[(2'h3):(2'h3)] >>> (-(8'hba)))) : ($signed($signed(wire60)) ?
              ({(8'h9c), (8'h9f)} ?
                  (wire67 ^~ wire62) : $signed(wire65)) : $signed($signed(wire65))))))
        begin
          reg73 <= $unsigned(wire57[(3'h7):(2'h2)]);
        end
      else
        begin
          reg73 <= $unsigned($signed(wire71[(1'h1):(1'h1)]));
          reg74 <= $signed((($unsigned($signed((8'had))) ?
              wire65[(2'h2):(2'h2)] : wire63[(2'h2):(1'h0)]) & (!((~^wire65) ?
              reg73[(1'h1):(1'h0)] : $unsigned((8'hbc))))));
          reg75 <= (8'hb8);
        end
      reg76 <= $signed($signed($unsigned(((wire72 ?
          wire69 : wire58) + {reg73}))));
      reg77 <= ({$unsigned(wire62[(4'hc):(3'h7)]),
          wire69[(1'h0):(1'h0)]} + reg74);
    end
  always
    @(posedge clk) begin
      reg78 <= ((reg76 << {wire69, wire60}) ^~ ((~{(|reg76),
          (|wire66)}) << $unsigned({((8'ha7) >= (8'hac))})));
    end
  assign wire79 = {(^~(+$signed($unsigned(wire63)))),
                      ((((|wire65) ?
                              $unsigned(wire61) : (&(8'hbc))) ^ ($signed(reg74) ?
                              reg75 : $unsigned(wire72))) ?
                          $unsigned((&wire61[(5'h10):(2'h3)])) : ($unsigned(reg75[(2'h3):(1'h0)]) ?
                              $unsigned((!reg73)) : wire71))};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module32  (y, clk, wire37, wire36, wire35, wire34, wire33);
  output wire [(32'hb1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire37;
  input wire [(3'h4):(1'h0)] wire36;
  input wire [(5'h13):(1'h0)] wire35;
  input wire signed [(4'ha):(1'h0)] wire34;
  input wire signed [(3'h6):(1'h0)] wire33;
  reg signed [(5'h15):(1'h0)] reg51 = (1'h0);
  reg signed [(4'he):(1'h0)] reg50 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg49 = (1'h0);
  reg [(4'he):(1'h0)] reg48 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg47 = (1'h0);
  reg [(5'h14):(1'h0)] reg46 = (1'h0);
  reg [(4'hf):(1'h0)] reg45 = (1'h0);
  reg [(4'h8):(1'h0)] reg44 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg43 = (1'h0);
  reg signed [(4'he):(1'h0)] reg42 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire41;
  wire signed [(3'h6):(1'h0)] wire40;
  wire [(3'h6):(1'h0)] wire39;
  wire signed [(4'hb):(1'h0)] wire38;
  assign y = {reg51,
                 reg50,
                 reg49,
                 reg48,
                 reg47,
                 reg46,
                 reg45,
                 reg44,
                 reg43,
                 reg42,
                 wire41,
                 wire40,
                 wire39,
                 wire38,
                 (1'h0)};
  assign wire38 = wire37;
  assign wire39 = wire33;
  assign wire40 = (((~&{(+wire34), (wire37 || wire39)}) ?
                          ($signed((+wire35)) << $signed(wire35)) : wire33) ?
                      wire37 : (wire37[(4'h9):(4'h9)] || {$unsigned((~&wire38)),
                          $unsigned($unsigned(wire36))}));
  assign wire41 = (-$signed($unsigned(wire33[(1'h0):(1'h0)])));
  always
    @(posedge clk) begin
      if ($unsigned({$unsigned(wire36),
          ($unsigned($unsigned((8'hab))) ?
              wire37 : ($unsigned(wire39) != $signed((8'hb3))))}))
        begin
          reg42 <= ($unsigned(wire36[(1'h1):(1'h1)]) ?
              ((((wire40 >> (8'ha7)) || (8'hbf)) ?
                  (~|$unsigned((7'h40))) : (wire39[(1'h0):(1'h0)] ?
                      wire36 : (wire40 ?
                          (8'h9f) : wire38))) >>> $signed(wire41)) : wire36[(2'h2):(1'h1)]);
          reg43 <= {(~^(wire40 ? wire39 : $signed(wire33[(2'h3):(1'h1)])))};
          reg44 <= (8'hb9);
          if ($signed(wire37))
            begin
              reg45 <= (|wire34);
            end
          else
            begin
              reg45 <= $unsigned((reg43[(4'h8):(3'h6)] ?
                  ((^{reg43, (8'hae)}) ?
                      $unsigned($signed(wire37)) : {$unsigned(wire33),
                          ((8'hb6) << reg44)}) : (reg45[(2'h2):(1'h1)] < wire35[(5'h11):(4'hb)])));
              reg46 <= {reg44[(3'h6):(1'h1)],
                  $unsigned({wire36, $signed(wire34[(1'h0):(1'h0)])})};
              reg47 <= (($signed($signed(wire41[(3'h5):(2'h2)])) ?
                  (~^wire40[(1'h1):(1'h0)]) : reg43) - (&wire35[(3'h5):(1'h1)]));
              reg48 <= {$unsigned($unsigned(wire37[(4'ha):(4'ha)])),
                  (({((8'ha9) ? wire36 : reg47), {(8'hb6), wire40}} ?
                          ((reg47 ? reg42 : wire33) ?
                              $signed(reg42) : $signed((8'hb3))) : wire37[(1'h0):(1'h0)]) ?
                      {({reg46, wire41} ?
                              reg44 : $signed(wire36))} : ({(wire38 >>> reg42)} - wire40[(3'h6):(2'h3)]))};
              reg49 <= reg44;
            end
        end
      else
        begin
          reg42 <= {(~&wire36), wire34[(3'h4):(3'h4)]};
          reg43 <= ((^~$signed((8'had))) | ($signed(((8'hb0) ~^ (reg47 & (8'hb2)))) <<< {wire34[(3'h4):(3'h4)],
              wire40}));
          reg44 <= ($signed(reg46) << $signed(wire37));
          if ($signed(($signed((~^$unsigned(reg47))) ~^ {$unsigned({reg45}),
              ((reg42 ~^ (8'hbd)) == reg43[(3'h6):(2'h3)])})))
            begin
              reg45 <= (-(~&wire38));
              reg46 <= (~&($signed((8'haf)) ^~ (~&((wire38 ?
                  wire40 : reg49) ~^ $signed(reg47)))));
              reg47 <= $unsigned((({(reg42 ? wire33 : reg42),
                  (~^wire37)} >>> (&wire35[(5'h10):(4'hc)])) < (wire36 ?
                  $signed(reg42) : $signed({reg49}))));
            end
          else
            begin
              reg45 <= $signed((reg48[(4'h9):(2'h2)] ?
                  (reg46[(4'h8):(1'h0)] ?
                      $signed(wire37) : ((reg45 ? reg42 : wire33) ?
                          reg49 : (+reg42))) : $signed($unsigned($unsigned(wire35)))));
              reg46 <= wire33[(3'h5):(2'h2)];
              reg47 <= $signed((reg49 <= (((reg44 ?
                  wire39 : reg42) > (|wire37)) ~^ reg48[(3'h7):(2'h3)])));
              reg48 <= $unsigned(reg44);
              reg49 <= wire35[(4'he):(4'ha)];
            end
        end
      reg50 <= $unsigned($signed(wire39[(3'h4):(3'h4)]));
      reg51 <= reg43[(3'h6):(2'h2)];
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module13
#( parameter param29 = (((({(8'hb8)} ? ((8'hb8) | (8'ha1)) : {(8'hbb)}) ~^ (((8'haa) ? (8'ha5) : (8'hbd)) ? ((8'hba) && (7'h40)) : ((8'hbe) ? (8'hb7) : (8'h9e)))) ? (&(((8'ha9) << (8'hb7)) ? ((8'hb1) <<< (8'h9e)) : (-(8'hba)))) : (^((&(8'hb2)) > ((8'hb3) * (8'hb8))))) ? (({((8'hbb) ? (8'hbe) : (8'hb7)), ((7'h43) ? (8'hbe) : (8'hb9))} ? (~|((8'hb2) & (8'hb6))) : (7'h41)) || ((((8'hb8) ? (8'ha7) : (8'ha7)) ? {(7'h42)} : ((8'haa) ? (8'hae) : (8'hb5))) & ({(8'ha4), (7'h42)} - ((8'hba) ? (7'h41) : (8'ha7))))) : (((!(+(8'hb3))) ? ((~^(7'h41)) || ((8'h9f) ? (8'hb8) : (8'hb6))) : (((8'ha8) * (7'h42)) ? {(8'ha5), (8'h9f)} : ((8'ha2) ~^ (8'hb2)))) >> ((((8'h9e) == (8'hb2)) != {(7'h44)}) ? (((8'ha7) ^~ (8'hb1)) >> ((8'hab) ? (8'ha6) : (8'haa))) : ((!(8'ha6)) - (8'hb3))))) )
(y, clk, wire17, wire16, wire15, wire14);
  output wire [(32'h76):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire17;
  input wire signed [(5'h13):(1'h0)] wire16;
  input wire signed [(4'hb):(1'h0)] wire15;
  input wire signed [(2'h3):(1'h0)] wire14;
  reg [(2'h3):(1'h0)] reg28 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg27 = (1'h0);
  reg [(4'hf):(1'h0)] reg26 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg25 = (1'h0);
  reg [(2'h3):(1'h0)] reg24 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire23;
  wire signed [(5'h12):(1'h0)] wire22;
  wire signed [(4'hd):(1'h0)] wire21;
  wire signed [(3'h4):(1'h0)] wire20;
  wire [(4'he):(1'h0)] wire19;
  wire signed [(4'he):(1'h0)] wire18;
  assign y = {reg28,
                 reg27,
                 reg26,
                 reg25,
                 reg24,
                 wire23,
                 wire22,
                 wire21,
                 wire20,
                 wire19,
                 wire18,
                 (1'h0)};
  assign wire18 = (({$unsigned(wire16[(4'hd):(4'hb)])} >> wire14[(1'h0):(1'h0)]) != $unsigned($unsigned((~^$signed(wire16)))));
  assign wire19 = $signed($unsigned(wire15));
  assign wire20 = $unsigned($unsigned(wire19[(4'ha):(3'h6)]));
  assign wire21 = $signed((~|wire18));
  assign wire22 = wire20[(1'h1):(1'h1)];
  assign wire23 = (wire19 >> {$signed(((~|wire19) && $signed(wire21))),
                      ((^wire22) ^ (8'h9c))});
  always
    @(posedge clk) begin
      reg24 <= (~(8'hbf));
      reg25 <= (^(((wire18[(3'h6):(3'h4)] ? $unsigned(wire18) : (~&wire17)) ?
              wire15[(3'h5):(2'h3)] : (&((8'hb1) <<< (8'hbb)))) ?
          ($unsigned($signed(wire18)) << ($signed(wire20) ?
              (wire14 ?
                  wire14 : wire20) : $signed((7'h42)))) : ((^~$signed((8'hab))) ?
              (+$unsigned(wire23)) : ((wire18 ? reg24 : wire19) ?
                  {(8'ha0), wire15} : wire15))));
      if (reg24)
        begin
          reg26 <= (~|($signed((wire21 && (!reg25))) && (!($signed(wire16) ?
              {(7'h41)} : (wire22 < wire16)))));
        end
      else
        begin
          reg26 <= ((-$unsigned({wire20, (^wire18)})) - (wire18 ?
              $signed((~(&wire21))) : (wire19[(4'h8):(3'h4)] ?
                  $unsigned($unsigned(wire22)) : (^((8'hb3) || (8'hac))))));
          reg27 <= wire18;
        end
      reg28 <= (|((wire19[(4'he):(2'h2)] ?
          wire16[(3'h6):(2'h3)] : ((+wire18) ^~ (wire23 ?
              wire17 : reg25))) != $signed(((!wire20) < (reg24 - wire16)))));
    end
endmodule