(* use_dsp48="no" *) (* use_dsp="no" *) module top
#( parameter param148 = ({(((8'hb0) != (8'hb6)) ? {{(8'hb5)}, (&(8'ha6))} : (~^(8'haa)))} >= ({{{(8'hb3)}, {(8'h9d)}}} * ((7'h41) <= {(~(8'h9d)), ((8'hb4) ? (8'hab) : (8'hac))})))
, parameter param149 = {((^(&((8'hbb) ? param148 : param148))) & ((8'hbe) >>> param148)), ({((param148 ? param148 : param148) == param148)} ? (8'ha1) : ((8'hb0) ? (param148 | (param148 ? (8'h9e) : (8'ha5))) : {{param148, param148}}))} )
(y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h1e0):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire4;
  input wire signed [(5'h10):(1'h0)] wire3;
  input wire [(5'h10):(1'h0)] wire2;
  input wire [(5'h13):(1'h0)] wire1;
  input wire signed [(4'ha):(1'h0)] wire0;
  wire [(2'h2):(1'h0)] wire147;
  reg [(4'hc):(1'h0)] reg146 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg145 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire98;
  wire signed [(5'h11):(1'h0)] wire6;
  wire signed [(4'hf):(1'h0)] wire5;
  wire signed [(5'h14):(1'h0)] wire100;
  reg signed [(5'h10):(1'h0)] reg101 = (1'h0);
  reg [(4'hf):(1'h0)] reg102 = (1'h0);
  reg [(3'h6):(1'h0)] reg103 = (1'h0);
  reg [(4'h8):(1'h0)] reg104 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg105 = (1'h0);
  reg [(5'h11):(1'h0)] reg106 = (1'h0);
  reg [(5'h10):(1'h0)] reg107 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg108 = (1'h0);
  reg [(4'he):(1'h0)] reg109 = (1'h0);
  reg [(4'h9):(1'h0)] reg110 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg111 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg112 = (1'h0);
  reg [(5'h13):(1'h0)] reg113 = (1'h0);
  reg [(5'h14):(1'h0)] reg114 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg115 = (1'h0);
  reg [(5'h12):(1'h0)] reg116 = (1'h0);
  reg [(4'hd):(1'h0)] reg117 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg118 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg119 = (1'h0);
  reg [(4'ha):(1'h0)] reg120 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg121 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg122 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg123 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg124 = (1'h0);
  reg [(4'hb):(1'h0)] reg125 = (1'h0);
  reg [(4'hf):(1'h0)] reg126 = (1'h0);
  reg [(5'h14):(1'h0)] reg127 = (1'h0);
  reg [(4'hf):(1'h0)] reg128 = (1'h0);
  wire [(2'h3):(1'h0)] wire143;
  assign y = {wire147,
                 reg146,
                 reg145,
                 wire98,
                 wire6,
                 wire5,
                 wire100,
                 reg101,
                 reg102,
                 reg103,
                 reg104,
                 reg105,
                 reg106,
                 reg107,
                 reg108,
                 reg109,
                 reg110,
                 reg111,
                 reg112,
                 reg113,
                 reg114,
                 reg115,
                 reg116,
                 reg117,
                 reg118,
                 reg119,
                 reg120,
                 reg121,
                 reg122,
                 reg123,
                 reg124,
                 reg125,
                 reg126,
                 reg127,
                 reg128,
                 wire143,
                 (1'h0)};
  assign wire5 = wire2;
  assign wire6 = (8'ha8);
  module7 modinst99 (wire98, clk, wire2, wire6, wire0, wire5, wire3);
  assign wire100 = (^~($signed($unsigned((8'h9d))) ?
                       (~((wire3 ? wire0 : wire4) ?
                           wire3[(4'he):(4'hd)] : (~wire3))) : (wire6[(4'hb):(3'h5)] ?
                           wire3 : ($signed(wire2) >= $unsigned(wire3)))));
  always
    @(posedge clk) begin
      reg101 <= (wire4 - $unsigned($signed((!(^wire6)))));
      if ({wire100[(5'h13):(1'h1)]})
        begin
          reg102 <= $unsigned($signed($unsigned(({wire98} ~^ (wire0 ?
              wire1 : wire3)))));
          reg103 <= reg101;
          reg104 <= $unsigned($unsigned(wire4[(2'h3):(1'h0)]));
          reg105 <= (^wire100);
        end
      else
        begin
          reg102 <= $signed($signed({wire100[(4'hb):(1'h1)],
              $unsigned($unsigned(wire6))}));
        end
      reg106 <= wire98;
    end
  always
    @(posedge clk) begin
      if ($unsigned({$signed((-wire5[(4'hb):(4'h9)])), (8'ha8)}))
        begin
          if (((wire100 <<< reg106[(3'h5):(1'h0)]) ?
              (($unsigned((wire6 ?
                      reg102 : (8'hae))) != reg101[(1'h1):(1'h1)]) ?
                  (&(((8'h9c) ?
                      wire4 : reg102) > (|wire2))) : $unsigned(reg101[(4'he):(3'h4)])) : (wire5 == $unsigned(reg101))))
            begin
              reg107 <= ((($unsigned($signed((8'ha0))) ?
                      (+(reg106 >>> reg105)) : (^~(wire98 ^ wire0))) <<< $unsigned((~&((7'h43) + wire6)))) ?
                  wire98[(4'hd):(4'h9)] : $unsigned((~(8'haf))));
              reg108 <= ($signed(reg103[(1'h0):(1'h0)]) + ($unsigned(reg106) > wire2));
              reg109 <= wire4[(1'h0):(1'h0)];
            end
          else
            begin
              reg107 <= $signed($unsigned((((wire3 ?
                      wire100 : wire1) & (reg107 <<< wire0)) ?
                  {wire3[(4'h9):(1'h0)],
                      $signed(wire2)} : reg104[(3'h4):(2'h3)])));
            end
          reg110 <= $signed($unsigned((((reg101 ? wire5 : wire0) ?
              wire1[(1'h0):(1'h0)] : (reg104 * reg101)) <= (^wire2[(4'hc):(4'h8)]))));
          if ((~&$unsigned($signed({$signed((8'hab)), {wire0, (8'ha9)}}))))
            begin
              reg111 <= ((^~(($unsigned(reg109) ?
                  reg104[(4'h8):(1'h1)] : (wire100 ?
                      reg110 : wire3)) ^~ (((7'h42) ~^ reg110) ?
                  $unsigned(reg108) : reg109[(3'h6):(2'h2)]))) * reg103[(1'h1):(1'h1)]);
              reg112 <= reg109[(3'h4):(1'h0)];
              reg113 <= ((({((8'hbe) < reg112),
                      (reg107 - (7'h41))} | $unsigned((^wire1))) && ($unsigned((wire1 ?
                      reg108 : wire98)) <= {(!(8'hab)), wire0})) ?
                  ($unsigned({(reg112 ? reg112 : wire100),
                      {wire100, wire6}}) >= wire4) : wire3[(4'hb):(2'h2)]);
              reg114 <= $signed(wire6);
            end
          else
            begin
              reg111 <= $signed($unsigned(wire1[(4'ha):(1'h0)]));
              reg112 <= $unsigned($signed((~|{reg110, $unsigned(wire6)})));
              reg113 <= $signed((reg101 + reg114));
              reg114 <= reg101;
              reg115 <= $unsigned((($unsigned((^~wire3)) << ((reg110 >= reg107) ?
                      (-reg103) : reg109)) ?
                  (reg102 ?
                      ((reg107 && wire4) ?
                          (reg112 ?
                              reg102 : wire98) : (reg105 && wire2)) : (-(+wire4))) : {$unsigned((~^wire5)),
                      (8'hb4)}));
            end
        end
      else
        begin
          reg107 <= $signed(reg104[(1'h0):(1'h0)]);
          if ((^~$signed(reg105[(2'h3):(1'h0)])))
            begin
              reg108 <= reg109;
            end
          else
            begin
              reg108 <= ($unsigned(reg105[(3'h7):(1'h0)]) - ($signed((~|(wire3 ?
                      reg115 : wire0))) ?
                  wire100 : ((wire1[(4'h8):(2'h2)] ?
                          ((7'h42) | reg115) : {reg107}) ?
                      ($unsigned(reg103) ?
                          (-reg104) : $signed(reg103)) : $unsigned($signed(wire1)))));
              reg109 <= (^~{$signed(reg110)});
            end
          reg110 <= (reg113 ?
              $unsigned(wire6) : {$unsigned($unsigned({wire98, (8'hbc)}))});
          reg111 <= $unsigned($signed((wire4[(1'h1):(1'h1)] ?
              reg113[(1'h0):(1'h0)] : wire0)));
          reg112 <= ($unsigned((({reg113, reg105} ?
                  $signed(reg113) : $unsigned(wire3)) ^~ wire1)) ?
              $unsigned((((reg102 >>> wire3) > (|reg114)) ?
                  (+reg106[(4'ha):(1'h0)]) : (~^wire3))) : wire6);
        end
      if (reg109)
        begin
          reg116 <= $signed(($signed((^~$unsigned((8'hb1)))) + reg112[(1'h1):(1'h1)]));
          if ((((reg107 != (reg107[(3'h4):(1'h0)] ?
                  (reg109 <= wire2) : reg109)) * (reg109[(2'h2):(2'h2)] ?
                  (reg109[(2'h3):(1'h1)] && (^reg109)) : reg112[(3'h5):(2'h2)])) ?
              reg116 : (^~{reg110, $unsigned((&wire2))})))
            begin
              reg117 <= {wire0[(2'h3):(2'h2)],
                  ($signed($unsigned(wire98)) ?
                      ((((8'hbd) >= wire100) ?
                          reg110 : (!reg102)) >= (-$signed(reg103))) : {{reg112[(3'h7):(3'h4)],
                              (reg109 >> reg109)},
                          wire5[(3'h5):(2'h2)]})};
            end
          else
            begin
              reg117 <= ((&(|reg105)) * reg102[(3'h6):(2'h2)]);
              reg118 <= reg104[(2'h2):(2'h2)];
              reg119 <= $signed(((wire6[(5'h10):(3'h7)] ?
                  (wire2 ?
                      $signed(wire0) : $unsigned((8'hb5))) : wire0) == ($unsigned(reg106[(1'h0):(1'h0)]) & $signed($unsigned(wire98)))));
            end
        end
      else
        begin
          if ((8'hbf))
            begin
              reg116 <= $unsigned(($signed(((reg108 ^ reg109) ?
                  (^~reg109) : (reg106 >= reg104))) << $unsigned(($signed(reg111) ?
                  (wire6 << wire4) : (wire1 < reg114)))));
              reg117 <= (($signed($signed(reg104[(3'h6):(3'h5)])) ^~ {(wire6[(4'he):(3'h5)] - (reg117 ^ (8'hbc)))}) ?
                  $unsigned((~$signed((!wire3)))) : (8'h9c));
            end
          else
            begin
              reg116 <= (~($unsigned(((reg109 + reg118) && (wire2 || wire0))) ?
                  reg109 : reg101[(4'hb):(1'h0)]));
              reg117 <= (!(wire4[(2'h3):(1'h1)] ?
                  {(wire3[(3'h6):(2'h2)] ?
                          reg102[(1'h1):(1'h0)] : $unsigned((8'ha3)))} : (!((reg117 ?
                      reg116 : wire1) == $unsigned(reg116)))));
              reg118 <= ((^$unsigned(reg104[(1'h0):(1'h0)])) >>> reg107[(3'h5):(1'h1)]);
              reg119 <= (&reg102);
            end
        end
      reg120 <= reg103;
      if (reg113[(1'h1):(1'h0)])
        begin
          reg121 <= ((reg113[(3'h4):(1'h1)] ?
              $unsigned((^~wire5[(3'h6):(2'h3)])) : reg120) <<< (((^reg105[(3'h7):(1'h0)]) != (^~(wire100 ?
                  reg109 : reg116))) ?
              ((&(reg105 ? reg108 : reg114)) ?
                  reg113[(2'h3):(2'h3)] : $unsigned(reg110)) : wire5));
          reg122 <= {wire98, {$signed({wire6[(3'h7):(2'h3)], (|wire1)})}};
          reg123 <= (8'hbd);
        end
      else
        begin
          if ((^$unsigned(reg107)))
            begin
              reg121 <= reg116[(3'h5):(2'h3)];
              reg122 <= (((reg120 << {$signed((8'ha2))}) ?
                      reg113 : (($unsigned(reg115) || (&reg109)) ?
                          reg114 : {(reg109 < wire3)})) ?
                  reg118[(3'h4):(2'h2)] : (+(^~(^{wire6, reg109}))));
              reg123 <= (wire0[(2'h2):(1'h0)] ~^ reg120);
              reg124 <= wire5[(4'h9):(4'h8)];
            end
          else
            begin
              reg121 <= (($signed(($unsigned(reg123) ? {(8'hb3)} : reg105)) ?
                  (^(reg114[(2'h3):(2'h2)] ?
                      reg120 : $signed(reg114))) : reg104[(4'h8):(1'h1)]) * reg111[(4'h8):(3'h6)]);
            end
          reg125 <= (!($signed(reg122[(4'hb):(2'h2)]) > reg113[(3'h5):(2'h3)]));
          reg126 <= (&(~$signed({$unsigned((8'hb0)), {wire1, wire6}})));
          reg127 <= (|(wire3[(4'hb):(2'h2)] ?
              $signed(({reg103, wire6} < reg125[(1'h1):(1'h1)])) : {{(~&reg126),
                      $signed(reg111)},
                  ({reg124} <= reg112)}));
        end
      reg128 <= $unsigned($unsigned(reg101[(4'hc):(4'hb)]));
    end
  module129 modinst144 (wire143, clk, reg102, reg106, reg127, reg107, reg113);
  always
    @(posedge clk) begin
      reg145 <= {wire4, (|wire5)};
      reg146 <= ($unsigned((reg145 << (reg103 < (reg121 ?
          (7'h42) : reg110)))) ^ reg106[(4'he):(2'h2)]);
    end
  assign wire147 = (~(((~|$signed(wire1)) ?
                           ((~|(8'hbd)) ~^ $unsigned(reg112)) : $unsigned($unsigned(reg118))) ?
                       {$unsigned((7'h42))} : $signed(wire2[(4'h8):(1'h0)])));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module129
#( parameter param142 = ((~((+(!(8'hbc))) ^~ (+((8'hbc) <= (8'hbd))))) ? {(({(8'hb5)} >>> ((8'hb9) ^ (8'ha4))) || ((-(8'ha2)) ? ((8'h9f) ? (8'had) : (8'hb9)) : ((7'h44) ? (8'ha0) : (8'ha3)))), ((((8'hb3) ? (8'hb9) : (8'haf)) != ((8'h9f) ? (8'hb0) : (8'ha9))) ? (~^(+(8'hbb))) : {((8'hb8) >> (8'hb4))})} : (~^(&(~&((8'hbd) * (8'hbb)))))) )
(y, clk, wire134, wire133, wire132, wire131, wire130);
  output wire [(32'h57):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h4):(1'h0)] wire134;
  input wire [(5'h11):(1'h0)] wire133;
  input wire [(5'h14):(1'h0)] wire132;
  input wire signed [(3'h5):(1'h0)] wire131;
  input wire [(5'h13):(1'h0)] wire130;
  wire signed [(5'h14):(1'h0)] wire141;
  wire signed [(3'h4):(1'h0)] wire140;
  reg [(5'h11):(1'h0)] reg139 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg138 = (1'h0);
  reg [(4'ha):(1'h0)] reg137 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg136 = (1'h0);
  wire [(4'h9):(1'h0)] wire135;
  assign y = {wire141,
                 wire140,
                 reg139,
                 reg138,
                 reg137,
                 reg136,
                 wire135,
                 (1'h0)};
  assign wire135 = ((8'hbd) >= (~&($signed((wire133 ?
                       wire133 : wire132)) > wire132)));
  always
    @(posedge clk) begin
      if (wire134[(1'h1):(1'h0)])
        begin
          reg136 <= wire132[(4'hf):(4'hb)];
          reg137 <= $signed((~wire131[(3'h4):(3'h4)]));
        end
      else
        begin
          reg136 <= wire134[(1'h1):(1'h1)];
        end
      reg138 <= (~|($signed(((wire134 ? reg137 : wire135) ?
          reg136 : (|wire134))) ^~ (((wire131 ?
          wire130 : wire130) <= (reg137 == wire131)) << $unsigned((-reg136)))));
      reg139 <= $unsigned({{$unsigned(((8'hb7) + wire135))}, wire133});
    end
  assign wire140 = wire134[(1'h1):(1'h0)];
  assign wire141 = (wire131[(3'h5):(1'h0)] ?
                       wire132[(5'h14):(4'hb)] : wire130[(1'h0):(1'h0)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module7
#( parameter param96 = (|({(((8'ha2) ? (8'hba) : (8'ha4)) ? (-(8'hbf)) : ((8'hbc) < (8'hb4)))} <= (8'haa)))
, parameter param97 = (~({({param96, param96} >>> param96), (^{param96, param96})} > {((param96 ? param96 : param96) - param96)})) )
(y, clk, wire12, wire11, wire10, wire9, wire8);
  output wire [(32'hd3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hc):(1'h0)] wire12;
  input wire signed [(5'h11):(1'h0)] wire11;
  input wire signed [(4'ha):(1'h0)] wire10;
  input wire signed [(4'hf):(1'h0)] wire9;
  input wire [(4'hf):(1'h0)] wire8;
  wire signed [(3'h4):(1'h0)] wire95;
  wire signed [(5'h12):(1'h0)] wire94;
  reg [(4'hc):(1'h0)] reg93 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg92 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg91 = (1'h0);
  reg [(5'h11):(1'h0)] reg90 = (1'h0);
  reg [(4'hf):(1'h0)] reg89 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg88 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg87 = (1'h0);
  reg [(5'h14):(1'h0)] reg86 = (1'h0);
  reg [(5'h10):(1'h0)] reg85 = (1'h0);
  reg [(2'h3):(1'h0)] reg84 = (1'h0);
  wire [(4'hc):(1'h0)] wire82;
  wire [(3'h5):(1'h0)] wire15;
  wire signed [(4'hb):(1'h0)] wire14;
  wire [(5'h15):(1'h0)] wire13;
  assign y = {wire95,
                 wire94,
                 reg93,
                 reg92,
                 reg91,
                 reg90,
                 reg89,
                 reg88,
                 reg87,
                 reg86,
                 reg85,
                 reg84,
                 wire82,
                 wire15,
                 wire14,
                 wire13,
                 (1'h0)};
  assign wire13 = $signed(wire10);
  assign wire14 = (+wire12);
  assign wire15 = $unsigned($signed({(^(!wire12))}));
  module16 modinst83 (wire82, clk, wire14, wire15, wire12, wire8);
  always
    @(posedge clk) begin
      reg84 <= (-wire10);
      reg85 <= ($signed($unsigned((+$unsigned((8'hbf))))) ^ $unsigned($signed((+((8'hb6) ?
          wire15 : wire11)))));
      if (wire82)
        begin
          reg86 <= (~&$unsigned(($signed({wire9}) ?
              wire9[(2'h2):(1'h1)] : {(8'hbf), $unsigned(wire14)})));
          reg87 <= {$unsigned({wire14[(3'h7):(3'h5)],
                  $unsigned((wire9 ? wire14 : wire10))}),
              ($signed(((reg84 ? (8'ha9) : reg85) ~^ $signed(wire10))) ?
                  ((~$signed(wire9)) ^ $signed({wire11})) : ($unsigned(wire15) ?
                      (&$signed(wire82)) : (8'h9d)))};
          if ((-(((~|wire14[(1'h0):(1'h0)]) ?
                  ($signed(wire13) ^ ((8'hb0) ? wire10 : wire8)) : reg87) ?
              $signed($signed((~|wire13))) : {(~wire10[(3'h7):(3'h5)]),
                  ((reg87 ? (7'h41) : (8'ha8)) ~^ $unsigned(wire9))})))
            begin
              reg88 <= $unsigned($signed((|($unsigned(wire14) ?
                  {(8'hab)} : (wire14 ? (8'hb5) : (8'ha5))))));
              reg89 <= $signed($unsigned(wire11[(1'h0):(1'h0)]));
              reg90 <= (((wire11[(2'h2):(1'h0)] ^~ $unsigned(((8'hae) <<< wire14))) ?
                      wire9 : wire11[(5'h11):(5'h11)]) ?
                  (^~$unsigned($signed($unsigned((7'h40))))) : $signed({(&wire8[(4'hc):(4'hb)])}));
              reg91 <= wire12;
            end
          else
            begin
              reg88 <= {reg87};
              reg89 <= ({{(reg86 ~^ reg91), wire12[(3'h6):(2'h3)]},
                  ((wire11 ? (reg89 ? wire15 : reg85) : reg86) ?
                      $signed((reg91 >>> wire8)) : wire11)} && $unsigned($signed($signed({wire10,
                  reg91}))));
            end
        end
      else
        begin
          reg86 <= (reg89[(3'h5):(1'h1)] ?
              $signed($unsigned((&(wire8 ? wire14 : wire11)))) : (reg85 ?
                  ((reg89 ? reg90 : (7'h44)) + reg91) : {((wire14 >> reg84) ?
                          {wire13, reg84} : (wire82 <<< (8'hab)))}));
          reg87 <= (^(|reg91[(3'h5):(3'h4)]));
        end
      reg92 <= $unsigned($signed($unsigned(reg84[(1'h0):(1'h0)])));
      reg93 <= wire82[(1'h0):(1'h0)];
    end
  assign wire94 = (reg85 > $unsigned($signed($unsigned((reg85 ?
                      wire13 : wire11)))));
  assign wire95 = $unsigned({(|$signed(wire94)),
                      $signed(reg88[(2'h3):(1'h0)])});
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module16
#( parameter param81 = (!((^~((+(8'haf)) ? (7'h42) : (~|(8'ha2)))) <= ((8'haa) ? (((8'hb9) * (8'hb0)) ? {(8'hb5), (8'hb1)} : (~|(8'ha9))) : {(^~(8'ha4)), (&(8'hb0))}))) )
(y, clk, wire20, wire19, wire18, wire17);
  output wire [(32'h29b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire20;
  input wire [(3'h5):(1'h0)] wire19;
  input wire signed [(3'h6):(1'h0)] wire18;
  input wire [(4'hf):(1'h0)] wire17;
  wire signed [(2'h3):(1'h0)] wire80;
  wire signed [(4'hd):(1'h0)] wire79;
  reg signed [(5'h14):(1'h0)] reg78 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg77 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg76 = (1'h0);
  reg [(4'he):(1'h0)] reg75 = (1'h0);
  reg [(3'h5):(1'h0)] reg74 = (1'h0);
  reg [(4'ha):(1'h0)] reg73 = (1'h0);
  reg [(4'h8):(1'h0)] reg72 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg71 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg70 = (1'h0);
  reg [(4'hb):(1'h0)] reg69 = (1'h0);
  reg [(5'h11):(1'h0)] reg68 = (1'h0);
  reg [(3'h5):(1'h0)] reg67 = (1'h0);
  reg [(5'h10):(1'h0)] reg66 = (1'h0);
  reg [(2'h3):(1'h0)] reg65 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg64 = (1'h0);
  reg [(2'h3):(1'h0)] reg63 = (1'h0);
  reg [(5'h10):(1'h0)] reg62 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg61 = (1'h0);
  reg [(4'hc):(1'h0)] reg60 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg59 = (1'h0);
  reg [(2'h3):(1'h0)] reg58 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg57 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg56 = (1'h0);
  reg [(4'hb):(1'h0)] reg55 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg54 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg53 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg52 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg51 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg50 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg49 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg48 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg47 = (1'h0);
  reg [(4'he):(1'h0)] reg46 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg45 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg44 = (1'h0);
  reg [(5'h10):(1'h0)] reg43 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg42 = (1'h0);
  reg [(5'h15):(1'h0)] reg41 = (1'h0);
  reg [(5'h11):(1'h0)] reg40 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg39 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg38 = (1'h0);
  reg [(4'h9):(1'h0)] reg37 = (1'h0);
  reg [(3'h5):(1'h0)] reg36 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg35 = (1'h0);
  reg [(3'h5):(1'h0)] reg34 = (1'h0);
  reg [(3'h7):(1'h0)] reg33 = (1'h0);
  reg [(2'h2):(1'h0)] reg32 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg31 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg30 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg29 = (1'h0);
  reg [(2'h2):(1'h0)] reg28 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg27 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg26 = (1'h0);
  reg [(4'hc):(1'h0)] reg25 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire24;
  wire signed [(4'hd):(1'h0)] wire23;
  wire [(3'h6):(1'h0)] wire22;
  wire [(4'hc):(1'h0)] wire21;
  assign y = {wire80,
                 wire79,
                 reg78,
                 reg77,
                 reg76,
                 reg75,
                 reg74,
                 reg73,
                 reg72,
                 reg71,
                 reg70,
                 reg69,
                 reg68,
                 reg67,
                 reg66,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 reg55,
                 reg54,
                 reg53,
                 reg52,
                 reg51,
                 reg50,
                 reg49,
                 reg48,
                 reg47,
                 reg46,
                 reg45,
                 reg44,
                 reg43,
                 reg42,
                 reg41,
                 reg40,
                 reg39,
                 reg38,
                 reg37,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 reg32,
                 reg31,
                 reg30,
                 reg29,
                 reg28,
                 reg27,
                 reg26,
                 reg25,
                 wire24,
                 wire23,
                 wire22,
                 wire21,
                 (1'h0)};
  assign wire21 = (wire18 ?
                      ({(((8'hab) ? wire17 : wire18) < wire17),
                          wire20} ^ (({wire17, wire20} ^ (wire20 * wire18)) ?
                          $signed((8'hb2)) : ({wire19, wire18} ?
                              (wire17 ? wire17 : wire19) : (wire19 ?
                                  wire20 : wire20)))) : $signed(wire17));
  assign wire22 = wire17;
  assign wire23 = wire22[(1'h0):(1'h0)];
  assign wire24 = (wire23 >= (8'had));
  always
    @(posedge clk) begin
      reg25 <= (~&((wire21[(4'h9):(4'h9)] <<< {{(7'h42), wire17},
          $unsigned((8'hb2))}) == (-wire17[(1'h0):(1'h0)])));
      if ($unsigned((!((!{(8'hb1)}) ?
          $signed($signed(wire24)) : ($unsigned(wire23) ?
              (-wire23) : wire23)))))
        begin
          reg26 <= (((wire17 * (~&$signed(wire24))) >> ((|(wire18 & (8'hbc))) ?
                  reg25 : {{wire19}})) ?
              (~^(~&(wire20[(4'h8):(3'h6)] >= $signed(wire18)))) : wire21);
          reg27 <= $signed((~|wire20[(3'h4):(1'h0)]));
        end
      else
        begin
          reg26 <= ($signed(wire17) ^ {((~(wire23 || wire17)) < {$signed(wire20),
                  (wire17 ~^ wire18)}),
              (7'h40)});
        end
      reg28 <= (^~$signed(wire23[(4'h9):(3'h6)]));
      reg29 <= (-$unsigned((^((7'h41) ?
          (wire17 && wire19) : (wire20 ? (7'h40) : (7'h42))))));
      reg30 <= ((^$signed(($unsigned(wire17) ?
              $unsigned(wire19) : (wire23 || wire19)))) ?
          (~wire24[(1'h0):(1'h0)]) : (^(~&{(&reg27), (&wire19)})));
    end
  always
    @(posedge clk) begin
      if ($unsigned($unsigned((!$unsigned($unsigned(reg28))))))
        begin
          reg31 <= ($signed((({reg26, reg30} ^ wire17[(1'h0):(1'h0)]) ?
              $unsigned($unsigned(reg29)) : wire24)) && (reg27[(3'h4):(2'h3)] | (^~reg26[(2'h2):(2'h2)])));
          reg32 <= ($signed((wire24 ?
                  $unsigned(wire20[(3'h6):(1'h1)]) : $signed($signed((8'h9e))))) ?
              {(~$signed(wire20))} : wire22[(1'h0):(1'h0)]);
          reg33 <= (^$unsigned($unsigned((reg28[(1'h1):(1'h0)] - $unsigned(wire19)))));
          reg34 <= reg25[(3'h7):(1'h0)];
          reg35 <= (reg26[(4'hf):(1'h0)] ^ $signed(wire23));
        end
      else
        begin
          reg31 <= {({({(8'ha6)} < $unsigned((8'hb2)))} >= wire21),
              reg31[(3'h5):(3'h4)]};
          reg32 <= $signed((({wire24[(2'h3):(2'h2)], (~wire23)} ?
              (((7'h42) == reg29) <<< reg26) : (~^{reg32, reg34})) == reg27));
          reg33 <= $signed((reg34[(1'h0):(1'h0)] * {((|reg27) * $signed(wire18)),
              ($unsigned(reg31) >>> reg33)}));
        end
      if ($signed(((~^($unsigned(wire19) != wire21[(2'h2):(1'h1)])) == wire20[(1'h0):(1'h0)])))
        begin
          reg36 <= (&((!($unsigned(reg28) | $unsigned(wire24))) != (wire20 != (8'haf))));
          reg37 <= wire21[(4'hc):(3'h7)];
          reg38 <= ($signed(reg25[(4'h9):(4'h9)]) || ($unsigned($unsigned(reg29[(1'h0):(1'h0)])) && ({{reg31,
                      wire17},
                  wire19} ?
              reg27[(2'h3):(1'h1)] : ((reg25 ? reg34 : wire23) ?
                  $signed(wire23) : (wire24 ? reg34 : (8'ha6))))));
          if ($unsigned($unsigned($signed($signed({reg34, reg30})))))
            begin
              reg39 <= reg30[(5'h10):(2'h3)];
              reg40 <= reg34;
              reg41 <= $unsigned($signed({reg26, reg28}));
              reg42 <= $unsigned(({$unsigned((^(8'h9c))),
                  ($signed(reg26) ?
                      wire19 : $unsigned(reg37))} - $unsigned($signed((reg27 > reg29)))));
            end
          else
            begin
              reg39 <= {((($unsigned(reg41) ?
                          $signed(reg25) : reg37[(4'h8):(1'h0)]) >>> ($signed(reg37) ?
                          (~&reg41) : (reg33 ? reg29 : reg28))) ?
                      reg26[(3'h5):(3'h5)] : (wire19 >>> ((reg36 ?
                          reg26 : reg39) ^ {reg33, reg32})))};
              reg40 <= $signed($unsigned({(reg33 >> (reg34 ? reg32 : reg25)),
                  wire19[(1'h0):(1'h0)]}));
              reg41 <= wire19;
              reg42 <= $unsigned((~^reg41[(4'ha):(1'h1)]));
            end
        end
      else
        begin
          reg36 <= ((reg28[(1'h0):(1'h0)] ?
              (|$signed(reg39[(1'h1):(1'h1)])) : $signed($signed(reg36))) > {reg28});
          reg37 <= wire24;
        end
      reg43 <= wire19;
    end
  always
    @(posedge clk) begin
      if (((-reg43[(4'h8):(4'h8)]) ~^ $unsigned(($signed((reg42 ?
          reg27 : (8'hb1))) >> ($signed(reg39) & (reg39 ~^ reg31))))))
        begin
          reg44 <= {reg39[(3'h6):(1'h1)], reg30};
          if ($signed({reg31,
              (reg32 ?
                  ($signed(reg27) ?
                      {wire19,
                          reg27} : $unsigned(reg33)) : $signed($unsigned((8'had))))}))
            begin
              reg45 <= (~$unsigned(((^~(reg43 ^~ wire19)) | ((~|reg28) ?
                  (+reg37) : (wire23 >> reg35)))));
              reg46 <= wire23[(2'h3):(1'h1)];
              reg47 <= (wire21 == (reg30[(5'h13):(2'h3)] ^~ wire24[(1'h0):(1'h0)]));
              reg48 <= reg45[(2'h3):(1'h0)];
            end
          else
            begin
              reg45 <= $unsigned(reg41);
            end
        end
      else
        begin
          if (({reg41, (reg42[(4'h8):(1'h0)] ^~ reg40)} ?
              reg44[(2'h2):(1'h0)] : (reg43 >>> reg38)))
            begin
              reg44 <= ($signed(($unsigned(((8'h9d) + wire24)) * ((&wire21) ?
                  $signed(reg45) : (8'ha8)))) * reg36[(1'h0):(1'h0)]);
              reg45 <= reg34;
            end
          else
            begin
              reg44 <= ($signed(((wire19 & (reg46 ? reg31 : (7'h43))) ?
                      (reg34 ?
                          reg34[(1'h1):(1'h0)] : reg35[(1'h0):(1'h0)]) : wire21)) ?
                  reg35[(5'h14):(3'h4)] : $unsigned($unsigned((^$signed(reg39)))));
              reg45 <= {reg48[(3'h4):(1'h1)],
                  (^~({$unsigned(reg34),
                      ((8'hb8) ? reg32 : reg46)} <= $signed($signed(wire19))))};
              reg46 <= (-reg32[(1'h0):(1'h0)]);
            end
          reg47 <= ((~&((~$signed(reg40)) ? wire24[(1'h0):(1'h0)] : wire24)) ?
              (|({(reg42 ? wire23 : reg36)} ?
                  $signed($signed(reg42)) : $unsigned($unsigned(reg33)))) : $signed({((reg34 ^~ wire23) * $unsigned(reg48)),
                  reg47[(3'h6):(3'h6)]}));
          if ((|reg27[(2'h3):(2'h3)]))
            begin
              reg48 <= reg48;
              reg49 <= (&(((|reg30[(3'h4):(1'h0)]) ?
                      {reg31[(4'h8):(2'h3)], {(8'h9e)}} : {(reg44 ?
                              wire19 : wire21)}) ?
                  wire20[(4'hb):(4'h8)] : {reg33}));
              reg50 <= (^(8'hac));
              reg51 <= ($unsigned((reg48[(4'ha):(4'h8)] - ($unsigned(reg45) ?
                  $signed(reg33) : $signed(reg36)))) < $signed(reg49[(4'h8):(3'h7)]));
              reg52 <= (wire17 ?
                  reg42 : $unsigned((wire22 ?
                      $unsigned((reg37 <<< reg48)) : ((^~(8'haa)) ?
                          $signed(reg34) : (reg25 ? (8'ha5) : reg29)))));
            end
          else
            begin
              reg48 <= {(($unsigned($unsigned(wire24)) ?
                          (~|(-reg26)) : {$signed((7'h42)),
                              (reg37 ^~ wire21)}) ?
                      ((reg40[(4'hc):(4'ha)] ?
                          $unsigned(reg41) : reg48) >= reg29) : $signed(((reg37 >= reg32) ?
                          (~reg38) : ((8'hb7) ? (7'h40) : wire19))))};
            end
        end
      reg53 <= $unsigned(((!$unsigned($unsigned(reg44))) ? reg46 : (~^reg31)));
      reg54 <= reg37;
    end
  always
    @(posedge clk) begin
      reg55 <= ($signed(reg49[(1'h1):(1'h1)]) ?
          reg36 : $unsigned({wire19,
              ($signed((8'hbd)) <<< (wire22 ? reg35 : reg40))}));
      reg56 <= reg42;
      reg57 <= (|wire21);
      if (reg43[(4'h8):(2'h2)])
        begin
          reg58 <= reg55[(3'h6):(1'h1)];
          reg59 <= ({((~^(reg52 >> reg36)) ?
                      (~|(!reg31)) : $signed((wire22 * reg28)))} ?
              {{(wire18 ~^ reg28)}} : (^~(~&reg55[(4'h9):(4'h9)])));
          if ({(^(reg41 ^~ (&$unsigned(reg51))))})
            begin
              reg60 <= ((-$signed({$unsigned(reg46), (reg41 <= reg51)})) ?
                  ($unsigned((|reg42)) != $unsigned((reg55 >= (!reg33)))) : ((|$unsigned($unsigned(reg30))) | (+wire18[(2'h2):(1'h1)])));
              reg61 <= $unsigned(reg42);
              reg62 <= ($signed((reg46 ?
                  $unsigned($unsigned(reg48)) : (reg49[(3'h4):(2'h3)] ^ (reg37 | reg46)))) ~^ reg55);
              reg63 <= $unsigned($unsigned(reg49[(1'h0):(1'h0)]));
            end
          else
            begin
              reg60 <= $signed(reg30);
            end
          reg64 <= reg55[(4'hb):(3'h5)];
          if (reg58[(1'h0):(1'h0)])
            begin
              reg65 <= (((reg42[(4'h9):(3'h7)] >> reg56[(1'h1):(1'h1)]) ?
                  $signed(($signed(wire17) ?
                      wire24 : reg40[(3'h4):(2'h3)])) : (-$unsigned((reg56 ?
                      reg44 : wire22)))) < (8'hbd));
              reg66 <= (wire19 ?
                  ((-reg54) >> ($signed({(8'ha5)}) ?
                      (((8'hb6) < (8'hbc)) <<< (reg51 ?
                          wire17 : (7'h41))) : ($unsigned(reg44) ?
                          $signed(reg26) : wire20[(4'h9):(4'h8)]))) : (reg43[(3'h6):(3'h5)] < {(&(8'ha2))}));
            end
          else
            begin
              reg65 <= (wire23[(1'h0):(1'h0)] != $signed((reg41 | {(-reg63)})));
              reg66 <= $signed(wire18[(2'h3):(1'h1)]);
              reg67 <= $signed({((reg35[(1'h1):(1'h1)] ?
                      ((8'hb4) ? wire23 : reg60) : {reg30,
                          reg50}) || reg47[(3'h7):(1'h0)])});
              reg68 <= reg59;
              reg69 <= (-($unsigned((reg67 ?
                  (!(8'ha5)) : reg44[(3'h4):(2'h3)])) >= (~&$signed($signed(wire20)))));
            end
        end
      else
        begin
          reg58 <= wire23;
          reg59 <= $unsigned(wire17);
        end
      if ((8'hb1))
        begin
          reg70 <= $signed(reg61);
          reg71 <= reg70[(1'h0):(1'h0)];
          reg72 <= $signed((8'ha3));
          if ((8'hae))
            begin
              reg73 <= ((reg33[(2'h3):(1'h0)] < reg61[(1'h0):(1'h0)]) ~^ ($unsigned($unsigned((reg29 ?
                  (8'hae) : reg39))) >>> reg59));
              reg74 <= (-$signed($signed((!$unsigned(reg58)))));
              reg75 <= (~^reg29);
              reg76 <= $signed(wire18[(3'h4):(2'h3)]);
              reg77 <= $signed(($unsigned((^$signed(wire20))) ?
                  reg27 : ($unsigned((reg53 ?
                      reg57 : reg28)) ~^ (!reg55[(4'hb):(2'h2)]))));
            end
          else
            begin
              reg73 <= (~|reg43[(5'h10):(1'h1)]);
            end
        end
      else
        begin
          reg70 <= ($signed((($signed(reg47) ^ (+reg58)) >> $unsigned((wire24 ?
              reg61 : (8'ha3))))) | (~&(($unsigned(reg50) >= ((8'hb5) ?
              (8'hbe) : reg57)) ^~ (-reg77[(4'hd):(4'h8)]))));
          reg71 <= (+$unsigned((reg60 <<< $unsigned(reg38[(3'h5):(1'h0)]))));
          reg72 <= ({(!(~&(reg73 ? wire17 : reg42))), reg71} ?
              ($signed((8'hac)) >>> $unsigned((reg45[(2'h3):(2'h3)] ?
                  $unsigned(reg27) : (reg60 ?
                      (8'hbf) : wire20)))) : (($signed((~&reg66)) ?
                  $unsigned(((8'ha7) == reg42)) : (-(reg65 ?
                      reg55 : wire19))) <<< (~^reg77)));
          if ((!reg53[(1'h1):(1'h0)]))
            begin
              reg73 <= $signed((reg62 ?
                  reg53 : ((~$signed(reg58)) ?
                      $signed((reg76 < reg30)) : {(|wire19),
                          $unsigned(reg27)})));
              reg74 <= $unsigned(reg48);
              reg75 <= $signed(reg71);
              reg76 <= $signed(reg63);
            end
          else
            begin
              reg73 <= {(8'hb7)};
              reg74 <= {$unsigned(reg72),
                  (~|(~&{reg75[(3'h7):(3'h5)], reg50}))};
              reg75 <= {reg58[(1'h0):(1'h0)], $signed((~(^~{reg77})))};
              reg76 <= {reg62};
              reg77 <= $unsigned($unsigned($unsigned((reg76 ?
                  (+reg47) : reg74[(1'h0):(1'h0)]))));
            end
          reg78 <= ((|$unsigned($unsigned($signed(reg46)))) << ((|{$signed(reg62)}) ?
              $signed((reg77 ?
                  reg42[(4'h8):(3'h6)] : $unsigned((8'ha4)))) : (reg69[(3'h6):(2'h2)] & $signed($signed(reg59)))));
        end
    end
  assign wire79 = reg31[(3'h7):(2'h3)];
  assign wire80 = ($unsigned((reg47[(3'h5):(2'h2)] || (-$signed(wire24)))) ?
                      ($signed($unsigned(reg56)) ?
                          ($unsigned((reg71 & reg51)) ?
                              ($signed(reg26) ^ wire18) : $signed(wire79[(2'h3):(2'h2)])) : (^{$signed(reg38)})) : (~^($unsigned($signed(reg34)) ~^ {reg25})));
endmodule