module top
#( parameter param484 = {({(8'hac), (((8'ha5) ? (8'hbb) : (8'haa)) ? (~^(8'hb0)) : ((8'hb0) - (8'hb9)))} ^~ (((8'hae) ? (~|(8'hbd)) : (~|(8'ha2))) ? (!((8'ha8) << (8'ha6))) : (((8'ha6) < (8'hb0)) ? (~(8'hac)) : (~^(8'had)))))}
, parameter param485 = (&param484) )
(y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h241):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hf):(1'h0)] wire3;
  input wire signed [(3'h4):(1'h0)] wire2;
  input wire [(5'h13):(1'h0)] wire1;
  input wire signed [(3'h5):(1'h0)] wire0;
  wire [(4'ha):(1'h0)] wire483;
  wire signed [(4'hb):(1'h0)] wire482;
  wire [(4'h9):(1'h0)] wire481;
  wire [(5'h11):(1'h0)] wire480;
  wire [(5'h15):(1'h0)] wire479;
  reg [(4'hc):(1'h0)] reg478 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg477 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg476 = (1'h0);
  reg [(5'h13):(1'h0)] forvar475 = (1'h0);
  reg [(3'h7):(1'h0)] reg474 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg473 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg472 = (1'h0);
  wire [(2'h2):(1'h0)] wire471;
  wire [(2'h2):(1'h0)] wire470;
  wire signed [(5'h13):(1'h0)] wire468;
  wire [(5'h13):(1'h0)] wire38;
  reg signed [(4'hd):(1'h0)] reg37 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg36 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg35 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg34 = (1'h0);
  reg [(5'h10):(1'h0)] reg33 = (1'h0);
  wire [(5'h13):(1'h0)] wire32;
  wire [(4'ha):(1'h0)] wire31;
  reg [(4'h9):(1'h0)] reg30 = (1'h0);
  reg [(2'h3):(1'h0)] reg29 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg28 = (1'h0);
  reg [(3'h7):(1'h0)] reg27 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg26 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire25;
  wire [(4'hd):(1'h0)] wire24;
  wire signed [(3'h5):(1'h0)] wire23;
  reg [(4'h9):(1'h0)] reg22 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg21 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg20 = (1'h0);
  reg [(4'ha):(1'h0)] reg19 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg18 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg17 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg16 = (1'h0);
  reg [(4'hc):(1'h0)] reg15 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar14 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg13 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar12 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg11 = (1'h0);
  reg [(4'ha):(1'h0)] forvar10 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg9 = (1'h0);
  reg [(3'h7):(1'h0)] reg8 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire7;
  reg signed [(5'h10):(1'h0)] reg6 = (1'h0);
  reg [(5'h11):(1'h0)] forvar5 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire4;
  assign y = {wire483,
                 wire482,
                 wire481,
                 wire480,
                 wire479,
                 reg478,
                 reg477,
                 reg476,
                 forvar475,
                 reg474,
                 reg473,
                 reg472,
                 wire471,
                 wire470,
                 wire468,
                 wire38,
                 reg37,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 wire32,
                 wire31,
                 reg30,
                 reg29,
                 reg28,
                 reg27,
                 reg26,
                 wire25,
                 wire24,
                 wire23,
                 reg22,
                 reg21,
                 reg20,
                 reg19,
                 reg18,
                 reg17,
                 reg16,
                 reg15,
                 forvar14,
                 reg13,
                 forvar12,
                 reg11,
                 forvar10,
                 reg9,
                 reg8,
                 wire7,
                 reg6,
                 forvar5,
                 wire4,
                 (1'h0)};
  assign wire4 = ($signed(({wire1[(4'hc):(4'h9)]} < wire2)) ?
                     $signed(wire3[(4'hb):(4'h8)]) : (^wire3));
  always
    @(posedge clk) begin
    end
  assign wire7 = reg6[(3'h5):(1'h0)];
  always
    @(posedge clk) begin
      reg8 = wire2;
      reg9 <= $unsigned($signed(wire3));
    end
  always
    @(posedge clk) begin
      for (forvar10 = (1'h0); (forvar10 < (3'h4)); forvar10 = (forvar10 + (1'h1)))
        begin
          reg11 <= (wire3 ?
              (forvar10[(4'h9):(1'h0)] ?
                  $signed(wire7[(2'h2):(1'h0)]) : {wire2[(1'h1):(1'h0)]}) : {$unsigned($unsigned($signed(reg6))),
                  $signed((&(wire7 ? wire4 : forvar5)))});
        end
      for (forvar12 = (1'h0); (forvar12 < (3'h4)); forvar12 = (forvar12 + (1'h1)))
        begin
          reg13 <= wire7[(2'h2):(2'h2)];
          for (forvar14 = (1'h0); (forvar14 < (2'h2)); forvar14 = (forvar14 + (1'h1)))
            begin
              reg15 <= $unsigned($signed(wire1[(3'h5):(3'h4)]));
              reg16 <= (({{forvar10}} ?
                  {forvar12,
                      (reg11 << reg11)} : ((forvar5[(4'h9):(4'h8)] > forvar5[(4'hb):(2'h2)]) ?
                      ($unsigned(wire0) & $unsigned(reg13)) : (wire4 == ((7'h41) > wire1)))) | $unsigned(reg11));
              reg17 <= reg8[(3'h4):(2'h2)];
              reg18 <= (~(wire3 + (8'hb0)));
              reg19 <= reg8[(3'h7):(1'h1)];
            end
          reg20 <= wire1[(1'h1):(1'h0)];
          reg21 <= (~|(!(8'hbf)));
        end
      reg22 <= reg17[(1'h0):(1'h0)];
    end
  assign wire23 = reg13[(4'h8):(2'h3)];
  assign wire24 = {{reg22[(2'h3):(2'h3)]},
                      (($unsigned((reg18 ? (8'h9f) : reg9)) ?
                              {(wire0 != reg19)} : reg20[(4'hd):(4'hc)]) ?
                          (8'h9d) : $unsigned(wire7[(2'h2):(2'h2)]))};
  assign wire25 = $unsigned(($signed($unsigned((reg13 <= reg13))) <= wire3[(3'h4):(1'h0)]));
  always
    @(posedge clk) begin
      reg26 <= (^($unsigned((-(reg8 <<< (7'h41)))) ^~ $signed(wire25[(3'h6):(1'h1)])));
      reg27 <= ((wire0[(1'h1):(1'h0)] ^ (reg13 | reg17[(1'h1):(1'h0)])) ?
          reg8 : (~(|(~^{wire4}))));
      reg28 <= (+reg8[(3'h6):(3'h6)]);
      reg29 <= (reg8[(3'h5):(3'h5)] > reg20);
      reg30 <= (^(reg15 ?
          $unsigned($signed(forvar12)) : (({wire2, forvar10} ?
                  $unsigned(reg28) : forvar14[(3'h6):(3'h4)]) ?
              {{reg17, wire7},
                  (wire0 * reg29)} : (wire23 << ((8'ha2) - wire2)))));
    end
  assign wire31 = wire1[(5'h11):(4'h8)];
  assign wire32 = ((^((|(wire0 * reg13)) < (wire23[(2'h3):(2'h3)] <<< $unsigned(reg17)))) ?
                      reg22 : $signed(reg9[(1'h0):(1'h0)]));
  always
    @(posedge clk) begin
      reg33 = (8'ha4);
      reg34 = {(&wire23),
          ($signed(((~|forvar14) ?
              $unsigned(reg11) : (reg18 ?
                  (8'hb8) : (8'hb2)))) <= ($unsigned($signed(reg19)) * $signed($signed(reg20))))};
      reg35 <= reg18[(3'h7):(3'h7)];
      reg36 <= (reg16 ?
          $signed({{$unsigned(reg6)}}) : (reg27 & $signed({(reg16 ?
                  reg17 : (8'h9c))})));
      reg37 <= reg30[(3'h7):(1'h1)];
    end
  assign wire38 = reg16[(3'h5):(2'h3)];
  module39 modinst469 (wire468, clk, forvar12, reg15, reg9, forvar10);
  assign wire470 = (^((((reg21 ? forvar5 : (8'hb7)) ?
                           (reg13 & reg30) : ((8'hb1) < wire23)) && (~|{wire2,
                           reg20})) ?
                       $unsigned($unsigned($signed(wire4))) : wire32[(4'he):(3'h7)]));
  assign wire471 = $unsigned($signed($unsigned((wire32 ? reg33 : reg33))));
  always
    @(posedge clk) begin
      reg472 <= reg17;
      reg473 <= $signed(reg26[(1'h1):(1'h1)]);
      reg474 <= reg19[(4'h9):(2'h2)];
      for (forvar475 = (1'h0); (forvar475 < (2'h2)); forvar475 = (forvar475 + (1'h1)))
        begin
          reg476 <= ($signed(reg30[(2'h3):(2'h3)]) >> ((~((reg11 ?
              (8'ha6) : (7'h41)) ^~ $signed((8'hb0)))) | $signed($signed($signed(wire32)))));
          reg477 = (reg13 + {reg473[(2'h2):(1'h0)]});
        end
      reg478 <= ($unsigned(reg19) ?
          (~&$unsigned($signed((^~reg6)))) : $signed((|reg15)));
    end
  assign wire479 = (~$unsigned($signed(wire0)));
  assign wire480 = ((wire479[(4'hd):(2'h2)] ?
                           ((forvar10 ?
                                   {forvar14, (8'hb4)} : (wire0 ?
                                       reg22 : reg17)) ?
                               wire24 : wire1) : reg37[(3'h7):(3'h4)]) ?
                       reg11 : (reg36[(2'h2):(1'h1)] ?
                           $unsigned(reg20[(4'hf):(4'h8)]) : $unsigned((|{wire7}))));
  assign wire481 = ($unsigned({reg20[(4'h9):(4'h8)],
                       ($signed((8'hbb)) ?
                           ((8'hb9) ?
                               reg20 : reg6) : (wire4 << reg473))}) <= (~|reg474[(1'h0):(1'h0)]));
  assign wire482 = (+reg36);
  assign wire483 = ((^~forvar5[(4'hd):(4'hd)]) >> forvar14[(5'h10):(3'h5)]);
endmodule

module module39
#( parameter param466 = (((({(8'ha1), (7'h42)} * (&(8'hb0))) ^~ (((8'ha8) < (8'hbb)) ? (8'haf) : ((8'ha6) << (8'h9d)))) || ((((7'h43) ~^ (7'h41)) ? ((8'haa) != (8'hb5)) : {(8'hba), (8'hb0)}) == ((&(8'hbd)) ? ((8'hab) <<< (8'hb9)) : (+(8'hb1))))) ? ((&({(8'h9f)} ? {(8'ha2), (8'ha3)} : ((8'hb4) ? (8'h9f) : (8'hbe)))) || ((~(^(8'haa))) > (((8'ha5) ? (8'hb6) : (8'h9d)) ? {(7'h40), (8'ha5)} : {(8'ha1)}))) : (~&{((~^(8'hb3)) ? (~(7'h42)) : (8'hbf)), {{(8'ha7)}, ((8'ha3) >>> (8'ha9))}}))
, parameter param467 = ({param466, (~^((param466 ? param466 : param466) << param466))} == (~&((~^((8'hb2) > param466)) ^~ ({param466, param466} == param466)))) )
(y, clk, wire40, wire41, wire42, wire43);
  output wire [(32'h33a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire40;
  input wire signed [(4'hc):(1'h0)] wire41;
  input wire [(3'h6):(1'h0)] wire42;
  input wire signed [(2'h3):(1'h0)] wire43;
  wire signed [(4'hd):(1'h0)] wire465;
  wire signed [(4'hb):(1'h0)] wire464;
  reg signed [(4'ha):(1'h0)] reg44 = (1'h0);
  reg [(3'h5):(1'h0)] reg45 = (1'h0);
  reg signed [(4'he):(1'h0)] reg46 = (1'h0);
  reg [(5'h11):(1'h0)] reg47 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg48 = (1'h0);
  reg [(5'h12):(1'h0)] reg49 = (1'h0);
  reg [(3'h4):(1'h0)] reg50 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire51;
  wire signed [(5'h14):(1'h0)] wire52;
  wire [(4'hd):(1'h0)] wire53;
  wire signed [(5'h15):(1'h0)] wire54;
  reg [(4'hf):(1'h0)] reg55 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg56 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar57 = (1'h0);
  reg [(5'h10):(1'h0)] forvar58 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg59 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg60 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar61 = (1'h0);
  reg [(5'h10):(1'h0)] reg62 = (1'h0);
  reg [(4'he):(1'h0)] reg63 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg64 = (1'h0);
  reg [(4'hd):(1'h0)] reg65 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg66 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg67 = (1'h0);
  reg signed [(4'he):(1'h0)] reg68 = (1'h0);
  reg [(2'h2):(1'h0)] reg69 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg70 = (1'h0);
  reg [(2'h2):(1'h0)] reg71 = (1'h0);
  reg [(5'h10):(1'h0)] reg72 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire73;
  wire [(5'h12):(1'h0)] wire74;
  wire signed [(4'h8):(1'h0)] wire75;
  reg [(5'h12):(1'h0)] forvar76 = (1'h0);
  reg [(5'h11):(1'h0)] reg77 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg78 = (1'h0);
  reg [(4'hf):(1'h0)] reg79 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg80 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg81 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg82 = (1'h0);
  reg [(4'hc):(1'h0)] reg83 = (1'h0);
  reg [(3'h7):(1'h0)] reg84 = (1'h0);
  reg [(5'h14):(1'h0)] reg85 = (1'h0);
  reg [(5'h13):(1'h0)] reg86 = (1'h0);
  reg [(4'h8):(1'h0)] reg87 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar88 = (1'h0);
  reg [(5'h12):(1'h0)] reg89 = (1'h0);
  reg [(5'h14):(1'h0)] reg90 = (1'h0);
  reg [(4'h8):(1'h0)] forvar91 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg92 = (1'h0);
  reg [(5'h10):(1'h0)] forvar93 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg94 = (1'h0);
  reg [(5'h15):(1'h0)] reg95 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg96 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg97 = (1'h0);
  reg [(4'ha):(1'h0)] reg98 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg99 = (1'h0);
  wire [(4'he):(1'h0)] wire462;
  assign y = {wire465,
                 wire464,
                 reg44,
                 reg45,
                 reg46,
                 reg47,
                 reg48,
                 reg49,
                 reg50,
                 wire51,
                 wire52,
                 wire53,
                 wire54,
                 reg55,
                 reg56,
                 forvar57,
                 forvar58,
                 reg59,
                 reg60,
                 forvar61,
                 reg62,
                 reg63,
                 reg64,
                 reg65,
                 reg66,
                 reg67,
                 reg68,
                 reg69,
                 reg70,
                 reg71,
                 reg72,
                 wire73,
                 wire74,
                 wire75,
                 forvar76,
                 reg77,
                 reg78,
                 reg79,
                 reg80,
                 reg81,
                 reg82,
                 reg83,
                 reg84,
                 reg85,
                 reg86,
                 reg87,
                 forvar88,
                 reg89,
                 reg90,
                 forvar91,
                 reg92,
                 forvar93,
                 reg94,
                 reg95,
                 reg96,
                 reg97,
                 reg98,
                 reg99,
                 wire462,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg44 <= (~^wire41[(1'h1):(1'h0)]);
      reg45 <= {{{{(~|reg44)}, ($unsigned(wire41) + $unsigned(wire42))},
              (!$unsigned((wire40 ~^ wire40)))},
          ($signed(wire40[(2'h2):(1'h1)]) ?
              (($unsigned(reg44) == ((8'ha9) ?
                  wire43 : wire43)) & wire43[(2'h3):(1'h0)]) : wire41)};
      reg46 <= wire41[(2'h2):(1'h0)];
      reg47 <= wire40;
    end
  always
    @(posedge clk) begin
      reg48 <= (+{$unsigned(($signed(reg45) ? (reg46 << reg45) : {reg44})),
          ($unsigned($unsigned(wire43)) ?
              ($unsigned(reg44) != $unsigned(wire42)) : (+(reg47 & reg47)))});
      reg49 <= wire40;
      reg50 = (^(|reg49[(2'h3):(1'h1)]));
    end
  assign wire51 = $unsigned({$signed(reg45[(3'h4):(3'h4)]),
                      ($signed($signed(reg48)) | {wire43})});
  assign wire52 = (|((|$signed($unsigned(wire51))) ^~ reg46));
  assign wire53 = reg47[(4'hd):(3'h7)];
  assign wire54 = (~^$unsigned($signed(reg48)));
  always
    @(posedge clk) begin
      reg55 <= (^~(^~($signed($signed(reg50)) >> (8'ha3))));
      reg56 = (((~|wire41[(3'h7):(3'h4)]) ?
          (8'hae) : (~|(~&$signed(wire51)))) * wire43);
      for (forvar57 = (1'h0); (forvar57 < (2'h3)); forvar57 = (forvar57 + (1'h1)))
        begin
          for (forvar58 = (1'h0); (forvar58 < (1'h0)); forvar58 = (forvar58 + (1'h1)))
            begin
              reg59 = $unsigned(wire41);
              reg60 <= forvar57;
            end
        end
      for (forvar61 = (1'h0); (forvar61 < (1'h1)); forvar61 = (forvar61 + (1'h1)))
        begin
          reg62 <= (|$unsigned(((reg55 ?
              (^~reg48) : wire42) >= (reg50[(1'h0):(1'h0)] >> $unsigned(reg49)))));
        end
    end
  always
    @(posedge clk) begin
      reg63 = $unsigned($signed(wire51[(4'hb):(1'h0)]));
      reg64 = (8'hbc);
      reg65 <= $unsigned({$unsigned((-$signed(forvar58)))});
      reg66 <= $unsigned(reg60[(2'h2):(1'h0)]);
      reg67 <= reg50[(1'h1):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg68 = (~|($unsigned((~^(forvar58 ?
          reg55 : reg48))) ^~ ((-(^forvar58)) >= (8'haf))));
      reg69 <= ($unsigned($signed({forvar57[(4'h8):(3'h5)], (~|(8'hb2))})) ?
          reg68[(3'h5):(3'h5)] : (reg44 ? (!reg67) : {(!(reg65 ~^ wire52))}));
      reg70 = $signed({(8'hb1), reg44[(3'h6):(2'h2)]});
      reg71 <= $unsigned($unsigned({($unsigned(reg62) ^ {wire51, reg59}),
          ({reg65, reg50} + {forvar58})}));
      reg72 <= (~&((((forvar58 ? (8'hbe) : reg46) * (forvar57 ?
                  reg68 : reg70)) ?
              ($unsigned(reg56) ? reg71 : $signed((8'ha0))) : {(~(8'hb7)),
                  $unsigned(reg60)}) ?
          ((8'hae) ?
              ((reg65 || reg66) ?
                  (reg69 ? reg55 : wire52) : (reg69 ?
                      reg50 : reg56)) : (+$signed(reg63))) : $signed(reg62[(3'h7):(3'h5)])));
    end
  assign wire73 = $signed(reg47[(1'h1):(1'h0)]);
  assign wire74 = reg62[(2'h3):(1'h0)];
  assign wire75 = ($unsigned(reg46[(4'he):(1'h0)]) != reg59[(1'h1):(1'h0)]);
  always
    @(posedge clk) begin
      for (forvar76 = (1'h0); (forvar76 < (3'h4)); forvar76 = (forvar76 + (1'h1)))
        begin
          if ((|($unsigned(wire51) ?
              $unsigned($signed((reg45 == wire73))) : ((^~(reg49 ?
                  wire52 : (8'ha9))) && {(reg46 * wire54)}))))
            begin
              reg77 <= $signed({($signed((wire43 ^ reg44)) <= (reg60[(4'hf):(2'h2)] ?
                      (reg60 >>> wire54) : {reg70}))});
              reg78 <= ((&{(+{wire42, reg69}), $signed((!reg70))}) ?
                  (reg46 < (((reg65 <<< wire40) - (+reg69)) >>> ((wire51 ?
                          (8'h9d) : forvar58) ?
                      (+forvar57) : reg60[(4'hc):(3'h5)]))) : (^$unsigned(reg59)));
              reg79 <= (~|($unsigned((|$unsigned(wire75))) | (8'ha9)));
            end
          else
            begin
              reg77 = ((&reg50) || wire54);
              reg78 <= (reg67[(1'h1):(1'h1)] != wire41);
              reg79 <= (~{$signed((^(reg71 ? reg50 : (8'hb9)))), wire43});
            end
          reg80 <= reg56[(3'h5):(1'h1)];
          if ((^(({(^reg68)} ?
                  (!$signed(wire42)) : (reg60[(1'h1):(1'h0)] && reg72)) ?
              {(((8'ha8) ? reg45 : forvar58) ?
                      (reg63 ? wire52 : reg71) : wire43),
                  {(reg50 ? (8'hbc) : reg68),
                      (wire53 ?
                          wire73 : reg77)}} : $unsigned(wire73[(4'ha):(3'h6)]))))
            begin
              reg81 = reg71;
              reg82 <= (reg68[(4'he):(4'he)] ?
                  ((^reg50) ?
                      reg71[(2'h2):(1'h1)] : ($signed(wire40) <<< (+reg81[(4'hd):(4'h9)]))) : (~(((reg65 <= wire43) <<< {reg67}) ?
                      {reg60} : (-((8'hbe) ? reg69 : (8'h9d))))));
              reg83 = (((~(wire51 << $signed((8'hb3)))) ?
                      ((reg47[(5'h10):(2'h3)] ?
                          $signed(reg70) : $signed(reg78)) != $unsigned((8'hb7))) : reg69) ?
                  reg66[(5'h11):(4'hf)] : {(reg48[(4'ha):(3'h5)] ?
                          (+reg47) : reg50)});
            end
          else
            begin
              reg81 = wire41;
            end
          reg84 <= {(!$unsigned((^~$unsigned(reg64))))};
          reg85 = reg45[(2'h2):(2'h2)];
        end
      reg86 = {$signed(wire43[(2'h3):(2'h3)])};
      reg87 <= reg66[(1'h1):(1'h0)];
      for (forvar88 = (1'h0); (forvar88 < (2'h3)); forvar88 = (forvar88 + (1'h1)))
        begin
          reg89 <= $unsigned(((7'h43) ?
              (((^wire73) ^ $signed(forvar88)) ?
                  ((reg80 != reg55) && $unsigned(wire54)) : (reg82 >>> $unsigned((7'h44)))) : $signed(((~&reg70) ?
                  $signed(reg77) : {(7'h40), wire54}))));
          reg90 <= $signed((^$unsigned(reg56)));
        end
      for (forvar91 = (1'h0); (forvar91 < (2'h3)); forvar91 = (forvar91 + (1'h1)))
        begin
          reg92 <= ({reg83[(3'h6):(2'h2)],
              (!($unsigned(reg77) + (reg70 ?
                  wire73 : wire53)))} & reg81[(4'hc):(2'h2)]);
        end
    end
  always
    @(posedge clk) begin
      for (forvar93 = (1'h0); (forvar93 < (2'h3)); forvar93 = (forvar93 + (1'h1)))
        begin
          reg94 <= (-(8'hba));
          reg95 = ((({$unsigned((8'ha1)), $signed(wire42)} ?
                      wire40 : (-$signed(reg55))) ?
                  ((8'hb8) ^~ ((reg83 ? reg48 : reg68) ?
                      {forvar61} : (~|wire43))) : $unsigned(((wire75 ?
                          reg85 : reg63) ?
                      (-reg80) : $signed(reg65)))) ?
              (forvar93 >= (~|(~forvar58[(4'h9):(4'h9)]))) : ((8'hbf) ?
                  (wire51[(4'ha):(3'h5)] <= reg67) : reg44[(3'h6):(2'h2)]));
          reg96 <= reg67;
          reg97 <= reg86[(3'h6):(2'h3)];
        end
      reg98 <= wire51[(4'hc):(3'h5)];
      reg99 <= {$unsigned(((^~((8'hae) ? wire51 : (7'h44))) == (^(reg64 ?
              reg67 : (8'hbc)))))};
    end
  module100 modinst463 (wire462, clk, forvar58, reg64, reg72, reg78, reg90);
  assign wire464 = ($signed($signed((8'hb3))) ^ wire74);
  assign wire465 = (8'hbf);
endmodule

module module100
#( parameter param461 = (!((|(((8'ha9) ? (8'hb3) : (8'hb2)) ? ((8'hb7) >> (8'hb0)) : {(7'h42)})) ? (!(&((8'hba) ? (8'hb0) : (8'hac)))) : ((~|(~(8'hbd))) ? (((8'hbb) ? (8'hbf) : (8'hba)) ? ((8'h9e) ? (8'hb9) : (8'hbd)) : ((8'ha0) ? (8'hae) : (8'h9e))) : (!((8'hab) ? (8'hb5) : (8'ha0)))))) )
(y, clk, wire101, wire102, wire103, wire104, wire105);
  output wire [(32'h2e9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire101;
  input wire signed [(2'h2):(1'h0)] wire102;
  input wire [(2'h2):(1'h0)] wire103;
  input wire signed [(5'h15):(1'h0)] wire104;
  input wire [(4'h8):(1'h0)] wire105;
  wire [(4'he):(1'h0)] wire460;
  wire signed [(4'h9):(1'h0)] wire459;
  wire [(4'hf):(1'h0)] wire458;
  reg [(2'h3):(1'h0)] reg457 = (1'h0);
  reg [(4'h8):(1'h0)] reg456 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg455 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg454 = (1'h0);
  reg [(5'h10):(1'h0)] reg453 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar452 = (1'h0);
  reg [(4'he):(1'h0)] reg451 = (1'h0);
  reg [(3'h6):(1'h0)] forvar450 = (1'h0);
  reg [(4'hf):(1'h0)] reg449 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire448;
  reg signed [(3'h5):(1'h0)] reg447 = (1'h0);
  reg signed [(4'he):(1'h0)] reg446 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg445 = (1'h0);
  reg [(5'h12):(1'h0)] reg444 = (1'h0);
  reg [(4'ha):(1'h0)] reg443 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg442 = (1'h0);
  reg [(5'h13):(1'h0)] reg441 = (1'h0);
  reg signed [(4'he):(1'h0)] reg440 = (1'h0);
  wire signed [(4'he):(1'h0)] wire439;
  wire signed [(4'hc):(1'h0)] wire106;
  wire signed [(4'h9):(1'h0)] wire107;
  reg [(4'hd):(1'h0)] reg108 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg109 = (1'h0);
  reg [(4'ha):(1'h0)] reg110 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg111 = (1'h0);
  wire [(5'h13):(1'h0)] wire112;
  reg signed [(5'h15):(1'h0)] forvar113 = (1'h0);
  reg [(4'ha):(1'h0)] reg114 = (1'h0);
  reg [(4'hb):(1'h0)] reg115 = (1'h0);
  reg [(3'h5):(1'h0)] reg116 = (1'h0);
  reg [(4'hc):(1'h0)] reg117 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg118 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg119 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg120 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg121 = (1'h0);
  reg [(3'h4):(1'h0)] reg122 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire123;
  reg signed [(4'h9):(1'h0)] reg124 = (1'h0);
  reg [(5'h10):(1'h0)] reg125 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg126 = (1'h0);
  reg [(4'ha):(1'h0)] reg127 = (1'h0);
  reg [(5'h13):(1'h0)] reg128 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar129 = (1'h0);
  reg [(5'h11):(1'h0)] reg130 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg131 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar132 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg133 = (1'h0);
  reg [(5'h12):(1'h0)] reg134 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg135 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg136 = (1'h0);
  reg [(3'h4):(1'h0)] reg137 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg138 = (1'h0);
  reg [(4'hc):(1'h0)] reg139 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg132 = (1'h0);
  reg [(5'h15):(1'h0)] reg140 = (1'h0);
  wire [(3'h7):(1'h0)] wire437;
  assign y = {wire460,
                 wire459,
                 wire458,
                 reg457,
                 reg456,
                 reg455,
                 reg454,
                 reg453,
                 forvar452,
                 reg451,
                 forvar450,
                 reg449,
                 wire448,
                 reg447,
                 reg446,
                 reg445,
                 reg444,
                 reg443,
                 reg442,
                 reg441,
                 reg440,
                 wire439,
                 wire106,
                 wire107,
                 reg108,
                 reg109,
                 reg110,
                 reg111,
                 wire112,
                 forvar113,
                 reg114,
                 reg115,
                 reg116,
                 reg117,
                 reg118,
                 reg119,
                 reg120,
                 reg121,
                 reg122,
                 wire123,
                 reg124,
                 reg125,
                 reg126,
                 reg127,
                 reg128,
                 forvar129,
                 reg130,
                 reg131,
                 forvar132,
                 reg133,
                 reg134,
                 reg135,
                 reg136,
                 reg137,
                 reg138,
                 reg139,
                 reg132,
                 reg140,
                 wire437,
                 (1'h0)};
  assign wire106 = $unsigned((8'haa));
  assign wire107 = (wire104[(4'hd):(3'h6)] >> (!(^$signed($signed((8'haa))))));
  always
    @(posedge clk) begin
      reg108 = (^$signed((~^$signed((wire102 ? wire102 : wire104)))));
      reg109 = {(~($unsigned({wire102}) && $unsigned($unsigned(wire105)))),
          ((wire106 <<< (&{(8'hb5)})) ^~ wire103)};
      reg110 <= $unsigned(($unsigned(wire101) ?
          (wire104 ^ ($signed(wire101) | $signed(wire105))) : ((~|$signed(wire106)) >= wire103)));
      reg111 <= wire104[(4'he):(1'h0)];
    end
  assign wire112 = (&{($unsigned(wire104[(4'hf):(1'h1)]) < (|((8'hb1) ?
                           reg110 : (8'ha8))))});
  always
    @(posedge clk) begin
      for (forvar113 = (1'h0); (forvar113 < (2'h2)); forvar113 = (forvar113 + (1'h1)))
        begin
          reg114 <= (($unsigned((&$unsigned(wire107))) ?
              wire102[(1'h0):(1'h0)] : $unsigned($unsigned((8'hbd)))) + (~&(((forvar113 | reg111) ?
              $signed(wire103) : (&(8'hba))) + reg110[(3'h6):(3'h5)])));
          reg115 <= ($unsigned((~^wire105)) ? reg114[(2'h2):(2'h2)] : wire107);
          reg116 <= $signed(reg109[(1'h0):(1'h0)]);
          reg117 <= (reg108 | $unsigned($unsigned(reg114)));
          reg118 <= $signed($signed(reg109[(3'h5):(1'h0)]));
        end
      reg119 <= (!reg117[(2'h3):(1'h0)]);
      reg120 <= $signed((((&(reg117 ?
          reg110 : (8'hb5))) - {(reg119 && (8'haf))}) >> $signed(($unsigned(reg109) ?
          $signed(reg114) : wire112))));
      reg121 <= ($signed(wire105[(3'h4):(2'h2)]) >> wire103[(2'h2):(1'h0)]);
      reg122 <= reg110[(3'h5):(3'h5)];
    end
  assign wire123 = (({$signed(reg110[(3'h4):(1'h1)]),
                               ((!reg116) < reg122[(3'h4):(2'h3)])} ?
                           ($unsigned(wire102[(1'h1):(1'h1)]) >= (^$signed((8'hb8)))) : (((!forvar113) + {wire107,
                               (8'hb2)}) <<< reg110)) ?
                       reg111[(2'h3):(2'h3)] : wire101[(3'h6):(1'h0)]);
  always
    @(posedge clk) begin
      reg124 <= $unsigned((({{reg120, reg117}} ?
              (~|$signed(wire123)) : ($signed(reg109) || $signed(reg110))) ?
          wire104 : reg115));
      reg125 <= $unsigned(wire123[(3'h6):(3'h4)]);
      reg126 <= wire123[(3'h4):(2'h3)];
    end
  always
    @(posedge clk) begin
      reg127 <= $unsigned((~&(+(reg117[(4'h9):(1'h0)] ?
          (8'ha6) : (reg116 | wire101)))));
      reg128 <= wire104;
      for (forvar129 = (1'h0); (forvar129 < (2'h2)); forvar129 = (forvar129 + (1'h1)))
        begin
          reg130 = reg121[(4'ha):(3'h6)];
          reg131 <= $signed((reg115 ?
              (((~|wire103) ?
                  (reg120 ?
                      reg130 : reg109) : ((7'h40) ~^ reg127)) <= {forvar129,
                  ((8'hb5) <<< wire103)}) : $unsigned((~|reg122[(1'h0):(1'h0)]))));
        end
      if (((wire106 ?
          ($signed(reg109[(3'h7):(3'h4)]) ?
              $signed(wire103) : $signed(reg130[(4'hf):(4'ha)])) : (((reg122 ~^ reg127) ?
                  $signed(reg120) : $unsigned((8'hb4))) ?
              (+(^forvar113)) : $signed((reg108 ?
                  reg115 : reg115)))) >>> $unsigned((($signed(wire123) > (^reg131)) >= $signed((wire102 ?
          wire106 : reg130))))))
        begin
          for (forvar132 = (1'h0); (forvar132 < (2'h3)); forvar132 = (forvar132 + (1'h1)))
            begin
              reg133 <= $unsigned({{{{forvar129, forvar113},
                          $signed(wire107)}}});
              reg134 <= reg109;
              reg135 <= (^~($signed(reg118[(4'h8):(1'h1)]) ?
                  (!{{wire101, reg115}, (wire102 < reg115)}) : reg133));
            end
          reg136 = ((~$signed(((wire106 ?
              reg131 : reg125) >= reg120))) + reg128);
          reg137 <= (wire103[(2'h2):(1'h1)] >> reg130[(4'he):(4'h8)]);
          reg138 <= ($signed({reg111[(1'h0):(1'h0)]}) ?
              $signed(($unsigned($signed(wire102)) ?
                  wire106[(1'h1):(1'h0)] : reg135[(1'h0):(1'h0)])) : reg115[(4'hb):(1'h1)]);
          reg139 <= reg122[(2'h2):(1'h0)];
        end
      else
        begin
          reg132 <= $signed($unsigned($signed((-$signed(reg114)))));
        end
    end
  always
    @(posedge clk) begin
      reg140 <= reg119;
    end
  module141 modinst438 (.wire144(wire104), .wire143(wire106), .wire145(reg135), .wire142(reg128), .clk(clk), .y(wire437), .wire146(wire112));
  assign wire439 = (~wire102);
  always
    @(posedge clk) begin
      reg440 <= reg111[(5'h12):(4'hb)];
      reg441 <= ($signed((reg120[(2'h3):(2'h2)] <= $unsigned((forvar132 ?
          forvar113 : reg108)))) && (($unsigned($signed(reg132)) != wire123) || reg127));
      reg442 <= $unsigned((|$signed($signed($signed((8'hbe))))));
      reg443 = forvar132;
    end
  always
    @(posedge clk) begin
      reg444 <= reg110[(3'h7):(2'h3)];
      reg445 <= {({forvar129} ?
              $unsigned($unsigned(reg134[(4'hf):(3'h6)])) : (reg444[(4'hf):(2'h2)] ?
                  wire106 : reg444[(4'hf):(4'ha)])),
          ($unsigned($signed($signed(reg440))) ?
              (&wire103) : ((&$unsigned(reg131)) - ($unsigned(reg128) <<< (~^reg125))))};
      reg446 <= $unsigned(reg120);
      reg447 <= ((~reg108) ^ (((((7'h41) << reg136) << (^wire105)) ?
              reg121 : $signed(wire102[(2'h2):(1'h0)])) ?
          reg110 : wire102[(1'h1):(1'h1)]));
    end
  assign wire448 = $signed($unsigned($unsigned($unsigned((&reg440)))));
  always
    @(posedge clk) begin
      reg449 <= $signed({$signed({{reg126}, $signed(reg447)}),
          {$unsigned({reg440})}});
      for (forvar450 = (1'h0); (forvar450 < (2'h3)); forvar450 = (forvar450 + (1'h1)))
        begin
          reg451 <= wire439;
          for (forvar452 = (1'h0); (forvar452 < (2'h3)); forvar452 = (forvar452 + (1'h1)))
            begin
              reg453 <= wire112;
            end
          reg454 <= reg126[(1'h1):(1'h1)];
          reg455 = (reg110 < ({reg126[(4'hb):(2'h3)],
              ((7'h43) != reg127)} - reg445[(4'hb):(3'h4)]));
          reg456 <= ((^((~&(8'had)) ?
                  $unsigned((reg134 ? (8'hbb) : reg131)) : $signed(reg134))) ?
              $signed($signed((8'h9d))) : reg134[(4'he):(2'h2)]);
        end
      reg457 <= $unsigned((&wire102));
    end
  assign wire458 = reg136;
  assign wire459 = $signed(reg441[(3'h6):(2'h3)]);
  assign wire460 = $unsigned((~^($signed(reg457) ?
                       reg111[(4'hb):(3'h5)] : $signed(reg125))));
endmodule

module module141
#( parameter param435 = ((^(((8'ha6) ? {(7'h41), (8'hb6)} : {(8'h9c), (8'hb7)}) ? {(&(8'h9d))} : {((8'h9f) ? (8'hbf) : (8'haf)), ((8'hb6) ? (8'hab) : (8'h9c))})) && ((~&(((8'hac) - (8'h9f)) ? ((8'ha1) ? (8'ha4) : (8'h9c)) : (^(8'hb8)))) ^ (+(8'ha9))))
, parameter param436 = (-(|(8'hab))) )
(y, clk, wire142, wire143, wire144, wire145, wire146);
  output wire [(32'h3f0):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h13):(1'h0)] wire142;
  input wire [(4'hc):(1'h0)] wire143;
  input wire signed [(4'hf):(1'h0)] wire144;
  input wire [(5'h14):(1'h0)] wire145;
  input wire signed [(5'h13):(1'h0)] wire146;
  wire [(4'ha):(1'h0)] wire434;
  reg signed [(3'h5):(1'h0)] reg433 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire432;
  reg signed [(3'h7):(1'h0)] reg431 = (1'h0);
  reg [(5'h10):(1'h0)] reg430 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg429 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg428 = (1'h0);
  reg [(3'h5):(1'h0)] reg427 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg426 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg425 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg424 = (1'h0);
  reg [(4'hd):(1'h0)] reg423 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg422 = (1'h0);
  reg [(3'h4):(1'h0)] reg421 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar420 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar419 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg418 = (1'h0);
  reg [(4'h8):(1'h0)] reg417 = (1'h0);
  reg [(4'h8):(1'h0)] reg416 = (1'h0);
  reg [(5'h11):(1'h0)] reg415 = (1'h0);
  reg [(2'h3):(1'h0)] reg414 = (1'h0);
  reg [(4'h9):(1'h0)] reg413 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar412 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg411 = (1'h0);
  reg [(4'hd):(1'h0)] reg410 = (1'h0);
  reg [(5'h10):(1'h0)] reg409 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg408 = (1'h0);
  reg [(4'hc):(1'h0)] reg407 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg406 = (1'h0);
  reg [(4'hf):(1'h0)] reg405 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar404 = (1'h0);
  reg [(4'hc):(1'h0)] reg403 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar402 = (1'h0);
  reg [(4'hc):(1'h0)] reg401 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg400 = (1'h0);
  reg [(3'h5):(1'h0)] reg399 = (1'h0);
  wire [(4'hc):(1'h0)] wire398;
  wire [(4'hd):(1'h0)] wire397;
  reg [(3'h6):(1'h0)] reg396 = (1'h0);
  reg [(2'h2):(1'h0)] reg392 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg395 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg394 = (1'h0);
  reg [(5'h11):(1'h0)] reg393 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar392 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg391 = (1'h0);
  reg [(5'h12):(1'h0)] reg390 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg389 = (1'h0);
  reg [(4'he):(1'h0)] reg388 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg387 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg386 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg385 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar384 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg383 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar382 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg381 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg380 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg379 = (1'h0);
  reg [(4'hf):(1'h0)] reg378 = (1'h0);
  reg [(4'he):(1'h0)] reg377 = (1'h0);
  reg [(5'h15):(1'h0)] forvar376 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg375 = (1'h0);
  reg [(4'hb):(1'h0)] reg374 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg373 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg372 = (1'h0);
  reg [(3'h4):(1'h0)] reg371 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg370 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar369 = (1'h0);
  reg [(5'h10):(1'h0)] reg368 = (1'h0);
  reg [(5'h10):(1'h0)] forvar367 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire147;
  wire [(4'hd):(1'h0)] wire148;
  reg [(5'h10):(1'h0)] forvar149 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg150 = (1'h0);
  reg signed [(4'he):(1'h0)] reg151 = (1'h0);
  wire [(5'h11):(1'h0)] wire152;
  wire [(2'h3):(1'h0)] wire153;
  reg [(5'h12):(1'h0)] reg154 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg155 = (1'h0);
  reg [(5'h10):(1'h0)] reg156 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire157;
  reg signed [(4'hc):(1'h0)] reg158 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg159 = (1'h0);
  reg [(5'h12):(1'h0)] reg160 = (1'h0);
  reg [(5'h15):(1'h0)] reg161 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg162 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg163 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg164 = (1'h0);
  wire [(4'h9):(1'h0)] wire365;
  assign y = {wire434,
                 reg433,
                 wire432,
                 reg431,
                 reg430,
                 reg429,
                 reg428,
                 reg427,
                 reg426,
                 reg425,
                 reg424,
                 reg423,
                 reg422,
                 reg421,
                 forvar420,
                 forvar419,
                 reg418,
                 reg417,
                 reg416,
                 reg415,
                 reg414,
                 reg413,
                 forvar412,
                 reg411,
                 reg410,
                 reg409,
                 reg408,
                 reg407,
                 reg406,
                 reg405,
                 forvar404,
                 reg403,
                 forvar402,
                 reg401,
                 reg400,
                 reg399,
                 wire398,
                 wire397,
                 reg396,
                 reg392,
                 reg395,
                 reg394,
                 reg393,
                 forvar392,
                 reg391,
                 reg390,
                 reg389,
                 reg388,
                 reg387,
                 reg386,
                 reg385,
                 forvar384,
                 reg383,
                 forvar382,
                 reg381,
                 reg380,
                 reg379,
                 reg378,
                 reg377,
                 forvar376,
                 reg375,
                 reg374,
                 reg373,
                 reg372,
                 reg371,
                 reg370,
                 forvar369,
                 reg368,
                 forvar367,
                 wire147,
                 wire148,
                 forvar149,
                 reg150,
                 reg151,
                 wire152,
                 wire153,
                 reg154,
                 reg155,
                 reg156,
                 wire157,
                 reg158,
                 reg159,
                 reg160,
                 reg161,
                 reg162,
                 reg163,
                 reg164,
                 wire365,
                 (1'h0)};
  assign wire147 = $unsigned($unsigned(((wire145 ^ wire144[(4'h9):(3'h4)]) << (^~(8'hb7)))));
  assign wire148 = (&$signed({{(wire146 + wire143)}}));
  always
    @(posedge clk) begin
      for (forvar149 = (1'h0); (forvar149 < (2'h2)); forvar149 = (forvar149 + (1'h1)))
        begin
          reg150 = (+wire145[(2'h3):(1'h1)]);
        end
    end
  always
    @(posedge clk) begin
      reg151 <= wire143;
    end
  assign wire152 = $signed(((!(~(forvar149 ? wire143 : wire143))) ~^ wire146));
  assign wire153 = (^({wire148[(4'hb):(3'h6)]} ?
                       $signed({$signed(reg151)}) : $signed((wire143[(4'h8):(3'h5)] - {wire148,
                           (8'hbb)}))));
  always
    @(posedge clk) begin
      reg154 <= ((!(+$signed(wire143[(3'h7):(2'h3)]))) > wire142[(5'h10):(1'h0)]);
      reg155 <= (($signed(reg154) >>> (-{wire144[(2'h3):(2'h2)]})) ?
          ($unsigned(((8'ha5) ?
              (~forvar149) : $signed(forvar149))) >>> wire153) : wire148);
      reg156 = (~^wire148[(4'hb):(3'h5)]);
    end
  assign wire157 = $unsigned(wire142);
  always
    @(posedge clk) begin
      reg158 = $unsigned($signed(((~^wire142[(2'h3):(1'h1)]) ^~ $signed($signed(reg155)))));
      reg159 <= ($signed(({(reg158 ? reg155 : wire153)} ?
              $unsigned((&reg151)) : $unsigned((reg155 >= reg154)))) ?
          ($signed((~^(!wire143))) < ((8'hb3) | $signed((&wire157)))) : wire153[(1'h0):(1'h0)]);
    end
  always
    @(posedge clk) begin
      reg160 = (~|wire145);
      reg161 <= (~|(wire143[(1'h0):(1'h0)] ?
          wire144 : ($signed($signed(wire143)) | $unsigned(reg159))));
      reg162 <= wire157[(4'h8):(3'h7)];
      reg163 <= ($unsigned((~reg151)) > $signed(reg156[(3'h7):(3'h5)]));
      reg164 <= (reg159[(4'hc):(4'hc)] != ($signed(((wire147 ?
              reg163 : wire152) << (reg160 <<< wire153))) ?
          $signed(reg163[(3'h5):(2'h2)]) : reg151[(4'hc):(4'h8)]));
    end
  module165 modinst366 (.wire167(reg151), .wire166(wire145), .wire170(reg158), .y(wire365), .wire169(wire148), .wire168(reg159), .clk(clk));
  always
    @(posedge clk) begin
      for (forvar367 = (1'h0); (forvar367 < (2'h3)); forvar367 = (forvar367 + (1'h1)))
        begin
          reg368 <= (reg163 ?
              reg163[(3'h6):(2'h2)] : $unsigned((&reg155[(4'ha):(3'h4)])));
        end
           for (forvar369 = (1'h0); (forvar369 < (1'h0)); forvar369 = (forvar369 + (1'h1)))
        begin
          reg370 <= $signed($signed(reg155));
          reg371 = reg158[(4'ha):(4'h9)];
          reg372 <= (~wire157[(4'h8):(2'h2)]);
          reg373 = (~^({(8'had)} != $signed((-(~|forvar369)))));
          reg374 <= reg158;
        end

    end
  always
    @(posedge clk) begin
      reg375 <= $signed(((forvar149 ? wire143 : (8'hab)) ?
          (+((wire147 - forvar369) < $signed(reg162))) : (^((wire365 * forvar367) ?
              reg372[(4'ha):(3'h6)] : (-wire143)))));
      for (forvar376 = (1'h0); (forvar376 < (2'h3)); forvar376 = (forvar376 + (1'h1)))
        begin
          reg377 <= ($signed({(^(forvar367 ?
                  wire142 : reg160))}) * (($unsigned((-reg372)) > $signed($unsigned(reg372))) + (+{{reg160,
                  reg159},
              {wire146}})));
          reg378 = ($signed((+({forvar367, reg375} ?
                  $unsigned(wire157) : reg163))) ?
              (reg375[(3'h7):(3'h7)] == reg158) : ({wire152,
                  reg368} <= {(~|$unsigned(wire145))}));
          reg379 <= reg368[(5'h10):(3'h4)];
        end
      reg380 <= reg374;
      reg381 <= $unsigned((~^(+reg370)));
      for (forvar382 = (1'h0); (forvar382 < (3'h4)); forvar382 = (forvar382 + (1'h1)))
        begin
          reg383 <= reg154[(1'h0):(1'h0)];
          for (forvar384 = (1'h0); (forvar384 < (1'h1)); forvar384 = (forvar384 + (1'h1)))
            begin
              reg385 <= (~&(reg156[(4'he):(2'h2)] > wire144[(1'h0):(1'h0)]));
              reg386 = $signed(((forvar369 + {wire144[(4'hd):(3'h6)],
                      (wire142 ? reg370 : (8'hbe))}) ?
                  ($signed(reg370[(4'hd):(1'h1)]) <<< (!reg370[(4'ha):(1'h1)])) : $signed(((reg385 && (7'h42)) ?
                      (wire157 <<< reg383) : (reg375 - reg158)))));
              reg387 = ($unsigned($signed($signed((~|reg150)))) == (forvar384 ?
                  reg374 : ($unsigned($signed(reg155)) ?
                      reg151[(1'h1):(1'h0)] : $signed((reg380 ?
                          reg378 : reg159)))));
              reg388 <= reg372[(4'ha):(2'h3)];
            end
          reg389 = ((|(-(forvar376 ? ((8'hbc) ^ reg380) : forvar369))) ?
              forvar382[(1'h1):(1'h0)] : (wire142 <= reg374));
        end
    end
  always
    @(posedge clk) begin
      reg390 <= reg383;
      reg391 <= forvar149;
      if ((~|($signed({$signed(reg389)}) <= $unsigned((8'hb2)))))
        begin
          reg395 = forvar384[(2'h3):(1'h1)];
        end
      else
        begin
          reg392 <= $signed(reg391[(1'h0):(1'h0)]);
          reg393 <= $unsigned(reg395);
          reg394 <= {{($signed(reg151) ?
                      $unsigned($unsigned(wire153)) : (+(reg393 ?
                          forvar392 : reg395)))},
              $signed((8'hb8))};
          reg395 <= $signed(reg373[(3'h4):(2'h2)]);
        end
      reg396 <= {reg151[(1'h1):(1'h0)],
          (-(reg374[(3'h5):(1'h0)] * ((reg163 > reg374) ^~ reg162[(3'h7):(2'h2)])))};
    end
  assign wire397 = $unsigned($signed($signed($unsigned((7'h40)))));
  assign wire398 = $unsigned(((~&$signed(wire152[(4'hc):(4'h8)])) ?
                       {$signed($unsigned((8'hb1))),
                           $unsigned(reg379[(1'h0):(1'h0)])} : $signed((+(reg390 ?
                           (8'hbd) : reg390)))));
  always
    @(posedge clk) begin
      reg399 <= {($unsigned((~&$unsigned(reg393))) ?
              ($unsigned(wire365[(2'h2):(2'h2)]) ?
                  ((reg377 != (8'hb1)) < reg159[(1'h0):(1'h0)]) : (~(wire365 != reg370))) : {reg391[(4'hd):(1'h0)]}),
          {(!$signed(reg372[(3'h6):(3'h6)])),
              ($unsigned(reg162[(3'h7):(3'h4)]) & $unsigned(reg389[(2'h3):(2'h3)]))}};
      reg400 <= wire153;
      reg401 <= ((-reg378[(4'hd):(3'h7)]) ?
          (8'ha3) : $signed((~$unsigned($unsigned((7'h42))))));
      for (forvar402 = (1'h0); (forvar402 < (2'h3)); forvar402 = (forvar402 + (1'h1)))
        begin
          reg403 <= ((reg383 ?
                  (reg155 ?
                      ((~^reg396) ~^ wire157[(3'h6):(1'h0)]) : $unsigned($unsigned(forvar149))) : wire145) ?
              (!({reg391,
                  (|reg391)} ^ (+wire397[(4'h8):(2'h2)]))) : $unsigned((reg391 > reg396[(2'h2):(2'h2)])));
          for (forvar404 = (1'h0); (forvar404 < (2'h3)); forvar404 = (forvar404 + (1'h1)))
            begin
              reg405 = reg370;
              reg406 <= reg374[(4'h9):(2'h2)];
              reg407 = (~(((((8'hb6) ? wire153 : wire142) == {reg161,
                      wire397}) >= $signed($unsigned(wire153))) ?
                  ({$unsigned(reg158)} ?
                      (8'ha5) : reg394[(2'h2):(1'h1)]) : (~$signed((8'ha6)))));
              reg408 <= ((!$signed($signed($unsigned((7'h40))))) > ($unsigned((8'h9d)) ?
                  {(-reg156[(4'ha):(3'h6)])} : {forvar392, reg388}));
            end
          reg409 <= $unsigned($unsigned(forvar367[(4'he):(3'h4)]));
          reg410 <= $unsigned((&(reg377[(4'ha):(4'h9)] ?
              ((forvar149 ? reg395 : (8'hbd)) >> $signed(reg393)) : {((8'hb2) ?
                      (8'hab) : wire147),
                  reg383[(4'hd):(4'hd)]})));
          reg411 <= {(reg389[(3'h4):(1'h1)] ?
                  (-forvar376[(5'h14):(4'he)]) : (~&$unsigned((reg156 ?
                      wire147 : reg403))))};
        end
      for (forvar412 = (1'h0); (forvar412 < (3'h4)); forvar412 = (forvar412 + (1'h1)))
        begin
          reg413 <= ($unsigned({($signed(reg399) ? (8'ha9) : (^~forvar402)),
                  reg374}) ?
              reg159[(3'h4):(2'h3)] : $signed($unsigned(reg394)));
          reg414 <= {$unsigned((^~forvar367[(3'h7):(1'h1)]))};
          reg415 <= reg380;
          reg416 <= reg371;
        end
    end
  always
    @(posedge clk) begin
      reg417 = {(reg394[(2'h2):(2'h2)] ?
              wire142 : ({$signed(wire144)} ?
                  (^(reg161 ? reg403 : reg393)) : wire398)),
          ((|$signed((wire145 ?
              (8'ha0) : reg411))) ~^ (((reg154 - reg151) ~^ (reg400 ?
              wire152 : reg163)) << $unsigned(reg394[(2'h2):(1'h0)])))};
    end
  always
    @(posedge clk) begin
      reg418 <= reg409;
      for (forvar419 = (1'h0); (forvar419 < (1'h1)); forvar419 = (forvar419 + (1'h1)))
        begin
          for (forvar420 = (1'h0); (forvar420 < (1'h0)); forvar420 = (forvar420 + (1'h1)))
            begin
              reg421 <= ((~|($signed({(8'hb7), wire147}) ?
                  $signed($unsigned(forvar404)) : reg408[(1'h1):(1'h1)])) - reg399[(2'h2):(1'h1)]);
              reg422 <= wire365;
              reg423 <= ((reg387 ? reg394 : reg151[(4'hd):(4'h8)]) ?
                  ({$signed((reg378 ? reg385 : reg164))} ?
                      {((-forvar149) * (forvar392 >> reg163))} : (((reg421 >> reg393) ?
                          $signed(reg417) : (reg374 ?
                              forvar420 : reg379)) ^ ((forvar376 + forvar420) <= (reg413 ?
                          reg164 : reg407)))) : (~&reg396[(2'h2):(2'h2)]));
              reg424 <= (~|reg160);
            end
          reg425 = ({(((reg370 * reg411) ? $signed(reg390) : $signed(reg158)) ?
                      $signed({reg383}) : wire142[(3'h5):(1'h1)]),
                  {(reg414 ~^ reg403), reg158}} ?
              $unsigned($unsigned($unsigned($unsigned(forvar382)))) : $signed(($unsigned({reg381,
                  reg424}) == $unsigned(((8'ha2) ? reg370 : wire153)))));
          reg426 = (+((((reg163 ? wire397 : wire365) - $unsigned(wire142)) ?
              wire153 : $signed((reg150 ?
                  reg423 : reg422))) >> forvar384[(3'h5):(2'h3)]));
          reg427 <= reg426[(1'h1):(1'h1)];
        end
      reg428 <= (wire157 != {(~reg372)});
      reg429 <= reg409;
      reg430 = $signed(reg390[(4'h9):(1'h1)]);
    end
  always
    @(posedge clk) begin
      reg431 = ((|reg421) > $signed(reg370));
    end
  assign wire432 = ($unsigned(forvar367) ?
                       $unsigned(reg430[(4'ha):(2'h3)]) : $unsigned((^(!$signed(reg408)))));
  always
    @(posedge clk) begin
      reg433 <= ($unsigned({$unsigned((8'hb0)),
          $signed((reg390 ^~ reg427))}) ^ $unsigned(($signed((reg392 < reg426)) ?
          reg156[(2'h2):(2'h2)] : (-(~^forvar384)))));
    end
  assign wire434 = (~^(reg406[(1'h1):(1'h0)] && reg163));
endmodule

module module165
#( parameter param363 = ((({{(8'hb7)}, (~&(8'ha9))} >= (!((8'hae) >> (8'h9d)))) || {({(8'ha8)} ? (8'h9c) : ((8'haf) + (8'hbc)))}) * {(((-(8'ha0)) ? (!(7'h43)) : (^~(8'hb1))) >> (^~{(8'hb8)})), {((-(7'h44)) > ((8'ha6) & (8'hbc))), (!((8'hbb) * (8'ha2)))}})
, parameter param364 = (&{param363}) )
(y, clk, wire170, wire169, wire168, wire167, wire166);
  output wire [(32'h298):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hc):(1'h0)] wire170;
  input wire signed [(4'hc):(1'h0)] wire169;
  input wire [(4'ha):(1'h0)] wire168;
  input wire signed [(4'hd):(1'h0)] wire167;
  input wire [(5'h14):(1'h0)] wire166;
  wire signed [(4'hf):(1'h0)] wire256;
  wire [(3'h6):(1'h0)] wire258;
  reg signed [(3'h6):(1'h0)] reg259 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg260 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg261 = (1'h0);
  reg [(3'h7):(1'h0)] reg262 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg263 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg264 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg265 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg266 = (1'h0);
  reg [(3'h6):(1'h0)] reg267 = (1'h0);
  reg [(3'h5):(1'h0)] reg268 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg269 = (1'h0);
  reg [(5'h14):(1'h0)] reg270 = (1'h0);
  reg [(5'h15):(1'h0)] reg271 = (1'h0);
  reg [(5'h14):(1'h0)] forvar272 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg273 = (1'h0);
  reg [(5'h10):(1'h0)] reg274 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire275;
  reg signed [(5'h14):(1'h0)] reg276 = (1'h0);
  reg [(4'hd):(1'h0)] reg277 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar278 = (1'h0);
  reg [(2'h3):(1'h0)] reg279 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg280 = (1'h0);
  reg [(3'h5):(1'h0)] reg281 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg282 = (1'h0);
  reg [(4'hc):(1'h0)] reg283 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg284 = (1'h0);
  reg [(3'h5):(1'h0)] reg285 = (1'h0);
  reg [(5'h11):(1'h0)] reg286 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg287 = (1'h0);
  wire [(4'h9):(1'h0)] wire288;
  reg signed [(3'h6):(1'h0)] reg289 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg290 = (1'h0);
  reg [(4'hd):(1'h0)] reg291 = (1'h0);
  wire [(5'h12):(1'h0)] wire292;
  reg signed [(5'h14):(1'h0)] forvar293 = (1'h0);
  reg [(5'h11):(1'h0)] reg294 = (1'h0);
  reg [(2'h3):(1'h0)] reg295 = (1'h0);
  reg [(5'h14):(1'h0)] reg296 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg297 = (1'h0);
  reg [(4'h9):(1'h0)] reg298 = (1'h0);
  reg [(5'h15):(1'h0)] reg299 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg300 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar301 = (1'h0);
  reg [(4'he):(1'h0)] reg302 = (1'h0);
  reg [(5'h14):(1'h0)] reg303 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar304 = (1'h0);
  reg [(4'he):(1'h0)] reg305 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg306 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg307 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg308 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg309 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar310 = (1'h0);
  reg [(2'h2):(1'h0)] reg311 = (1'h0);
  reg [(3'h5):(1'h0)] reg312 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire313;
  wire [(3'h6):(1'h0)] wire314;
  wire signed [(2'h3):(1'h0)] wire361;
  assign y = {wire256,
                 wire258,
                 reg259,
                 reg260,
                 reg261,
                 reg262,
                 reg263,
                 reg264,
                 reg265,
                 reg266,
                 reg267,
                 reg268,
                 reg269,
                 reg270,
                 reg271,
                 forvar272,
                 reg273,
                 reg274,
                 wire275,
                 reg276,
                 reg277,
                 forvar278,
                 reg279,
                 reg280,
                 reg281,
                 reg282,
                 reg283,
                 reg284,
                 reg285,
                 reg286,
                 reg287,
                 wire288,
                 reg289,
                 reg290,
                 reg291,
                 wire292,
                 forvar293,
                 reg294,
                 reg295,
                 reg296,
                 reg297,
                 reg298,
                 reg299,
                 reg300,
                 forvar301,
                 reg302,
                 reg303,
                 forvar304,
                 reg305,
                 reg306,
                 reg307,
                 reg308,
                 reg309,
                 forvar310,
                 reg311,
                 reg312,
                 wire313,
                 wire314,
                 wire361,
                 (1'h0)};
  module171 modinst257 (wire256, clk, wire169, wire166, wire170, wire168, wire167);
  assign wire258 = ($unsigned($signed(((wire256 ~^ (8'ha6)) ?
                           (wire166 != (8'hb4)) : (wire166 * (8'ha4))))) ?
                       {((~^(wire256 ? wire256 : wire167)) ?
                               {wire168[(3'h5):(3'h5)],
                                   (wire168 ? wire168 : wire168)} : (!{(8'hb3),
                                   wire168})),
                           ($unsigned((wire167 ?
                               wire256 : wire256)) >>> wire256[(4'h8):(4'h8)])} : $signed({(((8'hb1) ?
                                   wire168 : wire169) ?
                               $unsigned(wire169) : (~&wire169))}));
  always
    @(posedge clk) begin
      reg259 = (~|{(8'hbf)});
      reg260 = {({$unsigned($unsigned(wire167)),
              $signed((reg259 & wire168))} < ((-wire169[(3'h5):(3'h4)]) ?
              $signed((wire169 ? (8'hac) : reg259)) : $unsigned((-wire168)))),
          $signed(({$unsigned(wire258), wire168[(2'h3):(2'h2)]} ?
              (~^(~|(8'ha3))) : reg259[(3'h4):(3'h4)]))};
      reg261 <= wire170;
    end
  always
    @(posedge clk) begin
      reg262 = wire258[(1'h1):(1'h0)];
      reg263 <= $unsigned($unsigned($signed(wire170[(1'h0):(1'h0)])));
    end
  always
    @(posedge clk) begin
      reg264 <= wire168[(3'h5):(2'h2)];
      reg265 <= wire168[(4'h9):(4'h8)];
    end
  always
    @(posedge clk) begin
      reg266 = (reg263 ? reg263[(3'h7):(3'h6)] : (!$unsigned((8'ha3))));
      reg267 <= reg261;
      reg268 <= $signed(($signed(($signed(reg259) ?
          (wire169 ?
              reg261 : (8'hbc)) : (wire168 + wire170))) < ((+reg265[(3'h5):(2'h3)]) ?
          (~{wire258, wire167}) : {reg267[(2'h3):(2'h3)]})));
      reg269 <= ({((^~(~^reg264)) != (wire167 <= $signed(reg267))),
              (|(reg266[(3'h7):(2'h2)] * $unsigned(wire168)))} ?
          $unsigned($signed($signed($signed(reg263)))) : (-(8'ha0)));
    end
  always
    @(posedge clk) begin
      if (($signed(((reg265 ?
              {(8'ha0), reg264} : ((8'ha1) ? wire170 : (8'hb8))) ?
          (~wire166) : $signed($signed(reg265)))) <<< {(wire256[(4'hd):(2'h2)] & (wire167 ~^ (wire256 ~^ wire167))),
          {(~|(reg263 ? (8'h9e) : reg268))}}))
        begin
          reg270 <= (wire168[(1'h0):(1'h0)] ~^ ((wire166[(5'h10):(3'h7)] ?
                  $signed((reg268 || (8'ha2))) : (-(|(7'h42)))) ?
              (reg259 <<< $unsigned(reg269)) : (reg260[(2'h3):(1'h0)] | {(wire258 & reg263),
                  $signed((8'h9f))})));
          reg271 <= (|(|reg269[(4'hd):(1'h0)]));
        end
      else
        begin
          reg270 <= (|$signed((((reg266 ^ reg259) > wire167) < ($unsigned(reg264) ?
              wire166[(4'h9):(4'h9)] : (reg260 ? wire169 : reg262)))));
        end
      for (forvar272 = (1'h0); (forvar272 < (2'h2)); forvar272 = (forvar272 + (1'h1)))
        begin
          reg273 <= wire166;
        end
      reg274 <= $unsigned({$signed((^$signed(reg266)))});
    end
  assign wire275 = ((wire168 < ({reg268[(1'h1):(1'h1)]} ?
                           (reg263[(3'h6):(3'h4)] ?
                               reg265 : reg265) : $unsigned(reg270[(3'h6):(2'h2)]))) ?
                       ({reg261} ?
                           reg271 : reg269[(3'h4):(2'h3)]) : $signed($unsigned((8'haf))));
  always
    @(posedge clk) begin
      reg276 <= $signed(({(reg265[(3'h4):(2'h2)] == reg264),
          wire256} <<< $unsigned((|(wire166 ? reg273 : reg263)))));
      reg277 = (((~{(reg273 ?
              (8'h9c) : reg276)}) >>> wire167[(3'h6):(3'h6)]) || (8'hb9));
      for (forvar278 = (1'h0); (forvar278 < (2'h2)); forvar278 = (forvar278 + (1'h1)))
        begin
          reg279 <= (8'hbe);
          reg280 <= (8'ha0);
          reg281 <= (!$signed(((((8'ha2) ?
              wire275 : reg263) >> $unsigned(wire170)) | wire275)));
        end
      reg282 <= reg261;
      reg283 = $signed((&$signed(reg280)));
    end
  always
    @(posedge clk) begin
      reg284 = (7'h40);
      reg285 <= reg269;
      reg286 <= (|(~|($signed((&wire256)) ?
          ((reg279 <= reg266) ^~ $unsigned(reg269)) : $signed($unsigned((8'ha0))))));
      reg287 <= (8'ha5);
    end
  assign wire288 = forvar278;
  always
    @(posedge clk) begin
      reg289 = reg265[(3'h6):(3'h4)];
      reg290 <= $unsigned($signed($signed((~reg280))));
      reg291 = (8'hb2);
    end
  assign wire292 = (($unsigned({wire168[(1'h1):(1'h1)], (wire275 | reg265)}) ?
                           $signed((8'ha5)) : (~|$unsigned((wire258 ?
                               reg260 : reg268)))) ?
                       $unsigned((8'hb3)) : (((reg282 ?
                               reg271 : ((8'ha5) ^~ wire275)) ~^ reg269[(3'h5):(1'h1)]) ?
                           $signed(((8'hb3) ?
                               (reg285 * reg261) : (8'h9f))) : ($signed(wire167[(1'h1):(1'h1)]) ?
                               (&(^~wire258)) : (reg259 ?
                                   (reg286 ^ (8'ha2)) : (reg280 || reg263)))));
  always
    @(posedge clk) begin
      for (forvar293 = (1'h0); (forvar293 < (1'h0)); forvar293 = (forvar293 + (1'h1)))
        begin
          reg294 <= reg267;
          reg295 <= $signed((reg289[(3'h6):(3'h4)] <<< (reg273 ?
              $signed((+reg287)) : ((reg259 ? reg283 : reg259) ?
                  (reg266 <<< reg289) : $signed(wire167)))));
          reg296 = (reg281[(2'h2):(1'h0)] ? reg271 : $signed(reg264));
          reg297 = (($signed(reg273[(4'h8):(2'h3)]) ?
              (reg290 ?
                  ($signed(reg261) << {reg265, reg295}) : ({reg274, reg296} ?
                      (reg274 ?
                          wire169 : reg276) : (reg280 <<< reg262))) : (8'hbb)) - $unsigned($signed(($unsigned(reg266) && (wire168 ?
              reg282 : reg268)))));
        end
      reg298 <= ($unsigned(reg265) * {{reg285},
          $signed(((~(7'h43)) ? $unsigned(reg283) : {wire169}))});
    end
  always
    @(posedge clk) begin
      reg299 <= (wire256[(3'h7):(2'h3)] ?
          wire256 : ($signed((7'h43)) ?
              (((reg290 ? reg283 : (8'hb0)) ^ {reg297,
                  reg286}) == reg260) : ($signed($signed((8'ha3))) - ({wire275,
                      reg268} ?
                  {reg260} : $signed(reg286)))));
      reg300 <= reg286[(2'h3):(1'h0)];
      for (forvar301 = (1'h0); (forvar301 < (1'h0)); forvar301 = (forvar301 + (1'h1)))
        begin
          reg302 <= wire169;
          reg303 <= $signed((+{reg271, {(~^reg269), $signed((8'h9c))}}));
        end
      for (forvar304 = (1'h0); (forvar304 < (3'h4)); forvar304 = (forvar304 + (1'h1)))
        begin
          reg305 <= (forvar293 ? wire168 : $signed(reg290[(4'ha):(3'h5)]));
          reg306 <= $signed((~^reg285));
          reg307 <= (+(8'hb6));
        end
    end
  always
    @(posedge clk) begin
      reg308 <= (^~$signed($unsigned($signed({reg274}))));
      reg309 <= (reg290[(3'h6):(3'h4)] ?
          $signed($signed({$signed(reg262),
              (reg300 >= reg294)})) : $unsigned((^~{$unsigned(wire275)})));
      for (forvar310 = (1'h0); (forvar310 < (2'h2)); forvar310 = (forvar310 + (1'h1)))
        begin
          reg311 <= (($signed((~^$signed(reg266))) ?
              $unsigned({reg263, ((8'hb5) ? reg307 : reg279)}) : (~(reg299 ?
                  (&reg263) : reg271[(5'h13):(4'ha)]))) >>> {($unsigned((8'hbb)) ?
                  $signed((reg303 ?
                      wire168 : wire167)) : $signed($unsigned(forvar278))),
              reg270[(2'h3):(2'h3)]});
        end
      reg312 <= (reg276[(3'h4):(2'h3)] ?
          $signed((($signed(reg290) ? (reg308 && reg311) : $signed(wire292)) ?
              (~^{wire288, reg261}) : $unsigned((forvar293 ?
                  wire168 : wire258)))) : (!(~&$unsigned((reg284 ?
              reg298 : reg282)))));
    end
  assign wire313 = $signed(({(~&(~|reg283)),
                       $unsigned(reg305)} * (((&reg279) <<< $signed(reg306)) ?
                       {{reg260}, wire292} : (~^{reg289, reg270}))));
  assign wire314 = (!forvar272);
  module315 modinst362 (.wire319(reg273), .wire320(reg274), .clk(clk), .wire316(reg312), .wire317(reg259), .wire318(reg267), .y(wire361));
endmodule

module module315
#(parameter param360 = (8'hb7))
(y, clk, wire320, wire319, wire318, wire317, wire316);
  output wire [(32'h177):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire320;
  input wire [(4'hc):(1'h0)] wire319;
  input wire [(3'h6):(1'h0)] wire318;
  input wire signed [(3'h6):(1'h0)] wire317;
  input wire signed [(3'h4):(1'h0)] wire316;
  reg [(3'h6):(1'h0)] reg359 = (1'h0);
  reg [(4'hb):(1'h0)] reg358 = (1'h0);
  reg [(3'h7):(1'h0)] reg357 = (1'h0);
  reg [(4'he):(1'h0)] reg356 = (1'h0);
  reg [(3'h5):(1'h0)] reg355 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg354 = (1'h0);
  wire [(3'h7):(1'h0)] wire353;
  wire [(4'hb):(1'h0)] wire352;
  wire signed [(4'ha):(1'h0)] wire351;
  reg [(4'h9):(1'h0)] reg350 = (1'h0);
  reg [(4'hb):(1'h0)] reg349 = (1'h0);
  reg [(2'h3):(1'h0)] reg348 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg347 = (1'h0);
  reg [(5'h11):(1'h0)] reg346 = (1'h0);
  reg [(3'h4):(1'h0)] reg345 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg344 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg343 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg342 = (1'h0);
  reg [(2'h3):(1'h0)] reg341 = (1'h0);
  reg [(4'he):(1'h0)] reg340 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg339 = (1'h0);
  wire [(3'h6):(1'h0)] wire338;
  reg signed [(4'ha):(1'h0)] reg337 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg336 = (1'h0);
  reg signed [(4'he):(1'h0)] reg335 = (1'h0);
  reg [(2'h2):(1'h0)] reg334 = (1'h0);
  reg [(3'h5):(1'h0)] reg333 = (1'h0);
  reg [(4'ha):(1'h0)] reg332 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg331 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg330 = (1'h0);
  reg [(4'hb):(1'h0)] reg329 = (1'h0);
  reg [(4'hb):(1'h0)] forvar328 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg327 = (1'h0);
  reg signed [(4'he):(1'h0)] reg326 = (1'h0);
  reg [(5'h13):(1'h0)] forvar325 = (1'h0);
  reg [(4'hf):(1'h0)] reg324 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar323 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg322 = (1'h0);
  reg [(3'h5):(1'h0)] reg321 = (1'h0);
  assign y = {reg359,
                 reg358,
                 reg357,
                 reg356,
                 reg355,
                 reg354,
                 wire353,
                 wire352,
                 wire351,
                 reg350,
                 reg349,
                 reg348,
                 reg347,
                 reg346,
                 reg345,
                 reg344,
                 reg343,
                 reg342,
                 reg341,
                 reg340,
                 reg339,
                 wire338,
                 reg337,
                 reg336,
                 reg335,
                 reg334,
                 reg333,
                 reg332,
                 reg331,
                 reg330,
                 reg329,
                 forvar328,
                 reg327,
                 reg326,
                 forvar325,
                 reg324,
                 forvar323,
                 reg322,
                 reg321,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg321 = wire316[(2'h3):(1'h1)];
      reg322 = wire318;
      for (forvar323 = (1'h0); (forvar323 < (2'h2)); forvar323 = (forvar323 + (1'h1)))
        begin
          reg324 = (({($unsigned(wire316) ?
                          $unsigned(wire319) : (wire320 ? wire317 : wire318)),
                      wire319} ?
                  {wire316[(2'h2):(2'h2)]} : reg321[(2'h3):(1'h1)]) ?
              wire320[(4'hf):(4'hc)] : $unsigned(wire318));
        end
      for (forvar325 = (1'h0); (forvar325 < (1'h1)); forvar325 = (forvar325 + (1'h1)))
        begin
          reg326 <= wire319[(4'ha):(3'h5)];
          reg327 = (^~forvar323);
          for (forvar328 = (1'h0); (forvar328 < (1'h1)); forvar328 = (forvar328 + (1'h1)))
            begin
              reg329 <= wire317;
              reg330 = {forvar325};
              reg331 = (~&$signed(($unsigned((reg326 ?
                  forvar323 : wire317)) | ((!wire316) ?
                  ((8'h9d) << (8'ha0)) : {wire316}))));
            end
          reg332 <= $signed(wire316);
          reg333 <= (8'ha7);
        end
    end
  always
    @(posedge clk) begin
      reg334 <= forvar328[(1'h0):(1'h0)];
      reg335 = $unsigned({$signed({(reg324 << reg329)}),
          (wire316 ? (~{wire316, (8'hac)}) : (~$signed(forvar325)))});
      reg336 <= {($signed((8'hbf)) && reg331[(4'h8):(3'h6)]),
          reg335[(4'hb):(4'h9)]};
      reg337 <= reg332;
    end
  assign wire338 = $signed(reg332[(1'h1):(1'h1)]);
  always
    @(posedge clk) begin
      reg339 <= reg337;
      reg340 <= {reg330[(5'h10):(2'h3)]};
    end
  always
    @(posedge clk) begin
      reg341 <= $signed((~wire316[(2'h3):(2'h2)]));
      reg342 <= ($signed((({reg332, reg340} ?
                  reg332[(4'h8):(2'h2)] : (reg333 ? forvar323 : reg324)) ?
              ((wire319 <<< forvar328) > $unsigned((8'hb7))) : (~^$unsigned(wire320)))) ?
          (!((^(reg329 ? (8'hbb) : wire338)) ?
              {$unsigned(wire316),
                  (forvar328 ? reg334 : reg324)} : ((reg326 == wire317) ?
                  (-reg340) : forvar323[(5'h13):(5'h13)]))) : $signed(((8'ha0) ?
              $unsigned((reg337 < wire320)) : (|$unsigned(wire320)))));
      reg343 <= $unsigned(($unsigned(reg324[(4'h8):(4'h8)]) || wire318));
      reg344 <= $signed(wire320[(1'h1):(1'h1)]);
      reg345 <= (wire319[(1'h1):(1'h1)] ?
          $unsigned($signed((8'hbe))) : $signed((8'hb2)));
    end
  always
    @(posedge clk) begin
      reg346 <= wire316;
      reg347 <= wire338;
      reg348 <= (~$signed((($signed((8'hb4)) ?
          reg322[(4'h8):(2'h2)] : $unsigned(wire316)) & {wire338[(2'h2):(1'h1)],
          (~&reg329)})));
      reg349 <= (+((8'ha3) ?
          wire318[(2'h3):(1'h1)] : $signed(reg326[(3'h7):(3'h6)])));
      reg350 = {(wire320[(4'hc):(4'h9)] < reg330[(2'h2):(1'h1)]),
          reg322[(1'h0):(1'h0)]};
    end
  assign wire351 = (reg327 ? (~|reg333[(2'h3):(2'h3)]) : (8'hbc));
  assign wire352 = $signed(((~&wire338[(2'h3):(2'h3)]) ?
                       (~|reg336) : {$unsigned($unsigned((8'hb3))), reg327}));
  assign wire353 = reg335[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      reg354 = reg347;
    end
  always
    @(posedge clk) begin
      reg355 <= forvar323[(3'h6):(3'h4)];
      reg356 <= wire352[(4'h9):(2'h2)];
      reg357 <= $unsigned($signed((((!reg331) ?
          (~|reg349) : (7'h40)) ^~ $unsigned((wire316 ~^ reg334)))));
      reg358 = (((($unsigned((8'hb6)) ?
          {(8'hbf), (8'had)} : wire351) * wire351) <<< ((~^$unsigned(wire319)) ?
          (reg344[(3'h5):(1'h1)] | $signed(reg327)) : (!$signed((8'hbc))))) >> $unsigned(forvar323[(3'h7):(1'h1)]));
      reg359 <= reg324[(3'h7):(1'h0)];
    end
endmodule

module module171  (y, clk, wire176, wire175, wire174, wire173, wire172);
  output wire [(32'h379):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h2):(1'h0)] wire176;
  input wire signed [(5'h14):(1'h0)] wire175;
  input wire signed [(4'hc):(1'h0)] wire174;
  input wire [(3'h5):(1'h0)] wire173;
  input wire signed [(2'h3):(1'h0)] wire172;
  wire [(4'he):(1'h0)] wire255;
  wire [(5'h10):(1'h0)] wire254;
  reg signed [(4'h8):(1'h0)] reg253 = (1'h0);
  reg [(4'hb):(1'h0)] reg252 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg251 = (1'h0);
  reg signed [(4'he):(1'h0)] reg250 = (1'h0);
  reg [(5'h11):(1'h0)] reg249 = (1'h0);
  reg [(4'hb):(1'h0)] reg248 = (1'h0);
  reg [(2'h3):(1'h0)] reg247 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg246 = (1'h0);
  reg [(3'h5):(1'h0)] reg245 = (1'h0);
  reg [(3'h5):(1'h0)] reg244 = (1'h0);
  reg [(4'h8):(1'h0)] forvar243 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg242 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg241 = (1'h0);
  reg [(2'h2):(1'h0)] reg240 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg239 = (1'h0);
  reg signed [(4'he):(1'h0)] reg238 = (1'h0);
  reg [(4'h8):(1'h0)] forvar237 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar236 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg235 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg234 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar233 = (1'h0);
  wire [(4'hd):(1'h0)] wire232;
  wire [(4'hf):(1'h0)] wire231;
  reg signed [(2'h2):(1'h0)] reg230 = (1'h0);
  reg [(5'h14):(1'h0)] reg229 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg228 = (1'h0);
  wire [(2'h2):(1'h0)] wire227;
  reg signed [(5'h13):(1'h0)] reg226 = (1'h0);
  reg [(5'h10):(1'h0)] reg225 = (1'h0);
  reg [(5'h13):(1'h0)] reg224 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg223 = (1'h0);
  reg [(4'h9):(1'h0)] reg222 = (1'h0);
  reg [(5'h14):(1'h0)] reg221 = (1'h0);
  reg [(4'he):(1'h0)] reg220 = (1'h0);
  reg [(3'h5):(1'h0)] forvar219 = (1'h0);
  reg [(2'h2):(1'h0)] reg218 = (1'h0);
  reg [(2'h3):(1'h0)] reg217 = (1'h0);
  reg [(4'h9):(1'h0)] reg216 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar215 = (1'h0);
  reg [(2'h2):(1'h0)] forvar214 = (1'h0);
  reg signed [(4'he):(1'h0)] reg213 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar212 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg211 = (1'h0);
  reg [(4'hf):(1'h0)] reg210 = (1'h0);
  reg [(5'h11):(1'h0)] reg209 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg208 = (1'h0);
  reg [(4'hc):(1'h0)] forvar207 = (1'h0);
  reg [(5'h14):(1'h0)] forvar206 = (1'h0);
  reg [(5'h12):(1'h0)] reg205 = (1'h0);
  reg [(3'h4):(1'h0)] reg204 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg203 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg202 = (1'h0);
  reg [(4'h8):(1'h0)] reg201 = (1'h0);
  reg [(2'h3):(1'h0)] reg200 = (1'h0);
  reg [(2'h2):(1'h0)] reg199 = (1'h0);
  reg [(3'h6):(1'h0)] reg198 = (1'h0);
  reg [(5'h11):(1'h0)] forvar197 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar196 = (1'h0);
  wire [(5'h11):(1'h0)] wire195;
  wire signed [(5'h10):(1'h0)] wire194;
  reg [(3'h5):(1'h0)] reg193 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg192 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg191 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar190 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg189 = (1'h0);
  reg [(2'h2):(1'h0)] forvar188 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire187;
  reg [(4'hb):(1'h0)] reg186 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg185 = (1'h0);
  reg [(3'h6):(1'h0)] reg184 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg183 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire182;
  wire signed [(3'h5):(1'h0)] wire181;
  wire signed [(3'h4):(1'h0)] wire180;
  reg signed [(4'hb):(1'h0)] reg179 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg178 = (1'h0);
  wire [(4'hb):(1'h0)] wire177;
  assign y = {wire255,
                 wire254,
                 reg253,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 reg248,
                 reg247,
                 reg246,
                 reg245,
                 reg244,
                 forvar243,
                 reg242,
                 reg241,
                 reg240,
                 reg239,
                 reg238,
                 forvar237,
                 forvar236,
                 reg235,
                 reg234,
                 forvar233,
                 wire232,
                 wire231,
                 reg230,
                 reg229,
                 reg228,
                 wire227,
                 reg226,
                 reg225,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 forvar219,
                 reg218,
                 reg217,
                 reg216,
                 forvar215,
                 forvar214,
                 reg213,
                 forvar212,
                 reg211,
                 reg210,
                 reg209,
                 reg208,
                 forvar207,
                 forvar206,
                 reg205,
                 reg204,
                 reg203,
                 reg202,
                 reg201,
                 reg200,
                 reg199,
                 reg198,
                 forvar197,
                 forvar196,
                 wire195,
                 wire194,
                 reg193,
                 reg192,
                 reg191,
                 forvar190,
                 reg189,
                 forvar188,
                 wire187,
                 reg186,
                 reg185,
                 reg184,
                 reg183,
                 wire182,
                 wire181,
                 wire180,
                 reg179,
                 reg178,
                 wire177,
                 (1'h0)};
  assign wire177 = wire176[(2'h2):(1'h1)];
  always
    @(posedge clk) begin
      reg178 = ((~^wire172[(2'h3):(1'h1)]) ?
          ($unsigned({(wire176 * wire177), (wire174 << wire176)}) ?
              ($unsigned($unsigned(wire174)) > (((8'hb0) ? wire177 : wire174) ?
                  $signed(wire177) : (wire172 ?
                      wire174 : wire177))) : (($signed(wire173) ^ wire177[(4'h9):(3'h7)]) | wire176)) : wire175);
      reg179 = $signed((($signed(wire175) ?
              $unsigned(wire175) : ((+wire174) < reg178[(2'h3):(2'h2)])) ?
          $unsigned((!$signed(wire175))) : (wire172 > reg178[(3'h5):(2'h2)])));
    end
  assign wire180 = $signed(wire177);
  assign wire181 = $signed(wire173);
  assign wire182 = wire174;
  always
    @(posedge clk) begin
      reg183 = ($signed($unsigned($unsigned($signed(reg179)))) ^ wire176);
      reg184 <= wire176;
    end
  always
    @(posedge clk) begin
      reg185 = (~^(^$signed((reg183[(4'hc):(3'h5)] ?
          (reg183 != wire172) : reg184))));
      reg186 <= {$signed(reg185[(4'hb):(4'hb)])};
    end
  assign wire187 = ($signed((8'hb8)) ?
                       (~|(7'h41)) : {{$signed(wire182),
                               $signed(reg178[(2'h3):(1'h1)])}});
  always
    @(posedge clk) begin
      for (forvar188 = (1'h0); (forvar188 < (1'h1)); forvar188 = (forvar188 + (1'h1)))
        begin
          reg189 <= wire180[(1'h0):(1'h0)];
          for (forvar190 = (1'h0); (forvar190 < (2'h3)); forvar190 = (forvar190 + (1'h1)))
            begin
              reg191 = (wire174[(2'h3):(2'h3)] >> wire174);
              reg192 <= (+(wire174 ?
                  (~|(~^(-(8'hbd)))) : $unsigned(($signed(wire187) ?
                      $unsigned(wire175) : forvar190))));
              reg193 = wire182;
            end
        end
    end
  assign wire194 = (~&($unsigned($unsigned($signed(forvar190))) ?
                       ((forvar188 ?
                           (^~reg192) : $unsigned(wire176)) ~^ (8'ha3)) : $unsigned($signed(wire187[(1'h0):(1'h0)]))));
  assign wire195 = ($unsigned(wire181[(1'h0):(1'h0)]) ?
                       ($signed(reg183[(3'h6):(3'h5)]) ?
                           (reg192 ?
                               reg189[(3'h5):(3'h5)] : $signed($unsigned(reg191))) : ($signed($unsigned(wire175)) ?
                               {wire174} : (^wire180[(3'h4):(3'h4)]))) : (forvar190[(4'h8):(1'h1)] == ($signed((8'ha3)) >= $signed({wire182,
                           (8'hb6)}))));
  always
    @(posedge clk) begin
      for (forvar196 = (1'h0); (forvar196 < (1'h0)); forvar196 = (forvar196 + (1'h1)))
        begin
          for (forvar197 = (1'h0); (forvar197 < (2'h3)); forvar197 = (forvar197 + (1'h1)))
            begin
              reg198 = $unsigned(((7'h41) <<< (((wire174 ? reg184 : wire173) ?
                      (reg183 ^~ (8'ha0)) : wire174) ?
                  (8'hb4) : wire172)));
              reg199 <= reg185[(4'ha):(4'ha)];
              reg200 <= {($unsigned(wire195) ?
                      (($signed(reg191) >> (reg186 || wire181)) != reg183[(2'h2):(1'h0)]) : {$unsigned((reg193 ?
                              wire195 : (8'had))),
                          wire187})};
              reg201 = wire180[(2'h3):(2'h2)];
            end
          reg202 <= (-($signed((&$signed(wire180))) ? reg186 : (|reg198)));
          reg203 <= $signed($unsigned(((reg192[(3'h7):(3'h7)] >> $signed(wire182)) ~^ $signed((-reg183)))));
          reg204 <= ((forvar190 - wire177[(1'h0):(1'h0)]) ?
              {{({wire181} ? $signed((8'hb4)) : (&reg199)), {reg183}},
                  {($unsigned(reg202) ?
                          (wire180 ~^ reg185) : (wire187 ? wire175 : wire194)),
                      ($unsigned(wire175) ?
                          wire172 : $unsigned((8'hb1)))}} : (~(wire173[(2'h3):(1'h1)] ?
                  wire181[(3'h5):(1'h0)] : forvar197)));
          reg205 <= ($signed({$signed((wire194 ? reg193 : wire173))}) & reg179);
        end
      for (forvar206 = (1'h0); (forvar206 < (2'h3)); forvar206 = (forvar206 + (1'h1)))
        begin
          for (forvar207 = (1'h0); (forvar207 < (3'h4)); forvar207 = (forvar207 + (1'h1)))
            begin
              reg208 <= wire180[(3'h4):(1'h1)];
              reg209 <= reg185;
              reg210 <= ($unsigned((($unsigned(wire195) | reg178[(3'h7):(3'h6)]) == $signed($signed(forvar188)))) >>> ((8'ha4) - {wire174}));
              reg211 <= $unsigned({(reg208 ?
                      $signed((reg203 && reg189)) : reg199[(2'h2):(1'h1)]),
                  (~^$unsigned(wire175[(5'h13):(5'h13)]))});
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar212 = (1'h0); (forvar212 < (1'h1)); forvar212 = (forvar212 + (1'h1)))
        begin
          reg213 <= ($unsigned($signed((forvar190[(2'h3):(1'h1)] ?
                  (8'h9f) : $signed(reg211)))) ?
              {(^~((forvar212 ? (8'hbd) : (8'h9e)) ?
                      ((8'ha7) ? wire174 : reg203) : (reg210 ?
                          reg189 : forvar196)))} : (^$signed($unsigned($unsigned(reg202)))));
        end
      for (forvar214 = (1'h0); (forvar214 < (1'h1)); forvar214 = (forvar214 + (1'h1)))
        begin
          for (forvar215 = (1'h0); (forvar215 < (2'h3)); forvar215 = (forvar215 + (1'h1)))
            begin
              reg216 <= ((^$signed((!(forvar197 ? wire181 : forvar197)))) ?
                  $signed({reg210[(4'h8):(1'h0)]}) : ($signed(wire173[(1'h1):(1'h0)]) - $signed(reg183[(2'h2):(2'h2)])));
              reg217 <= reg185[(5'h12):(3'h5)];
            end
          reg218 = $unsigned($unsigned(forvar207[(4'hc):(3'h7)]));
          for (forvar219 = (1'h0); (forvar219 < (3'h4)); forvar219 = (forvar219 + (1'h1)))
            begin
              reg220 = $unsigned(((^{(reg216 | reg204)}) ?
                  wire175[(5'h14):(4'ha)] : wire194));
              reg221 = reg201;
              reg222 <= (^{$signed(wire175), forvar188});
            end
          reg223 <= reg222[(3'h7):(3'h7)];
        end
      reg224 <= reg213[(3'h7):(1'h0)];
      reg225 <= (reg210[(4'hf):(3'h4)] ?
          (((8'hb0) + $unsigned(reg186[(2'h2):(1'h0)])) | reg204[(2'h2):(1'h0)]) : (+$unsigned($signed(reg178))));
      reg226 <= wire195[(4'h9):(3'h6)];
    end
  assign wire227 = $unsigned(reg209);
  always
    @(posedge clk) begin
      if ((^$signed($unsigned($unsigned((^~wire176))))))
        begin
          reg228 <= ((wire177[(1'h0):(1'h0)] & reg217[(1'h1):(1'h1)]) > (~&{reg222,
              forvar215}));
          reg229 = wire172;
          reg230 = reg193[(2'h3):(1'h1)];
        end
      else
        begin
          reg228 <= ($signed($signed((~&(forvar212 | reg198)))) && (reg185 != reg223[(3'h6):(1'h0)]));
          reg229 <= $signed(reg201[(3'h5):(1'h0)]);
        end
    end
  assign wire231 = reg193;
  assign wire232 = ($unsigned((^~$signed((wire194 + reg218)))) + ((reg185 ?
                       $unsigned((wire227 ?
                           reg199 : forvar215)) : (~^$signed(reg185))) || ($unsigned($signed((8'hbc))) == $signed($signed(forvar196)))));
  always
    @(posedge clk) begin
      for (forvar233 = (1'h0); (forvar233 < (2'h3)); forvar233 = (forvar233 + (1'h1)))
        begin
          reg234 = $unsigned($signed((reg193[(3'h4):(1'h1)] ?
              $unsigned($unsigned(wire180)) : {(wire172 ? (8'hb1) : (8'h9f)),
                  reg218[(2'h2):(1'h1)]})));
          reg235 = ($unsigned(((|((8'ha2) && reg229)) > ((7'h41) == $signed((8'ha2))))) ^~ $unsigned($signed(reg184)));
        end
      for (forvar236 = (1'h0); (forvar236 < (1'h1)); forvar236 = (forvar236 + (1'h1)))
        begin
          for (forvar237 = (1'h0); (forvar237 < (3'h4)); forvar237 = (forvar237 + (1'h1)))
            begin
              reg238 <= ($unsigned((((~wire175) ?
                  wire175 : (reg200 ?
                      reg183 : reg199)) | $unsigned(reg211))) >= (-(wire194 ?
                  (&$signed(reg217)) : {reg204[(2'h2):(1'h0)]})));
            end
          reg239 = $unsigned(((8'hae) ~^ reg234[(4'h8):(1'h0)]));
          reg240 <= $unsigned((((forvar188[(1'h1):(1'h1)] ?
                      $unsigned(reg217) : wire174[(2'h3):(2'h2)]) ?
                  (wire187[(5'h10):(2'h3)] ?
                      (reg213 >>> wire177) : (reg208 ?
                          reg203 : reg198)) : (wire232 == reg189)) ?
              ((^{(8'h9d)}) ?
                  (~|(!reg229)) : $signed(reg210)) : $signed({(reg189 ?
                      reg184 : reg217),
                  ((8'h9f) <<< wire176)})));
          reg241 = (~|(!$unsigned((8'hb6))));
          reg242 = (|($unsigned($unsigned((+forvar188))) ^~ ($signed($unsigned(reg234)) >>> $signed($signed(reg192)))));
        end
      for (forvar243 = (1'h0); (forvar243 < (3'h4)); forvar243 = (forvar243 + (1'h1)))
        begin
          reg244 = $signed((((!reg189[(3'h4):(1'h0)]) ?
              (-(+reg183)) : ($signed(reg230) <= wire175[(4'h8):(3'h7)])) * $signed(reg184)));
        end
      reg245 = reg199[(1'h1):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg246 <= ((^~($unsigned(((8'hbd) ?
              reg229 : (8'ha8))) + (~&$unsigned(reg235)))) ?
          $signed(reg241) : $unsigned((^~$signed((~&reg178)))));
      reg247 <= $unsigned((!reg204));
      reg248 = wire175;
    end
  always
    @(posedge clk) begin
      reg249 <= {$signed((reg211[(4'hb):(2'h3)] ?
              $unsigned($unsigned(reg242)) : reg234))};
    end
  always
    @(posedge clk) begin
      reg250 = $signed(((~reg218[(2'h2):(1'h0)]) ?
          forvar214[(2'h2):(1'h1)] : $signed($unsigned($unsigned(reg208)))));
      reg251 = forvar212[(3'h7):(3'h5)];
      reg252 <= $signed(reg205);
      reg253 = {$unsigned($signed(((reg240 >>> (7'h44)) && (reg218 ~^ reg245)))),
          (~|(reg235[(4'hb):(3'h6)] && ((~reg178) <= reg216[(3'h5):(2'h2)])))};
    end
  assign wire254 = $signed(reg251[(4'hf):(4'hc)]);
  assign wire255 = forvar196[(4'h9):(3'h7)];
endmodule