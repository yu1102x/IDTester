(* use_dsp48="no" *) (* use_dsp="no" *) module top
#( parameter param462 = ({(|((!(8'hac)) << (-(7'h43))))} ? (~|(8'hab)) : {(({(8'hb4), (8'hbf)} > ((8'ha0) & (8'h9f))) ~^ (((8'hbb) < (8'ha4)) | (~|(7'h43)))), (^({(8'hb8)} << ((8'haf) ? (8'hbc) : (8'ha3))))})
, parameter param463 = ((|param462) ? ((|(^(param462 == (8'hb5)))) ? (param462 < ((~(8'ha2)) + (^param462))) : ((((8'h9f) * (8'h9e)) ? (param462 * param462) : param462) ? {((7'h42) ? param462 : param462)} : param462)) : param462) )
(y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h37c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h7):(1'h0)] wire3;
  input wire signed [(4'hf):(1'h0)] wire2;
  input wire [(4'h8):(1'h0)] wire1;
  input wire [(3'h7):(1'h0)] wire0;
  wire signed [(5'h14):(1'h0)] wire461;
  reg signed [(4'hf):(1'h0)] reg460 = (1'h0);
  reg [(4'ha):(1'h0)] reg459 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg458 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar457 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg456 = (1'h0);
  reg [(2'h2):(1'h0)] reg455 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar454 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg453 = (1'h0);
  reg [(4'hd):(1'h0)] reg452 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire450;
  reg [(4'hb):(1'h0)] reg71 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg70 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg69 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar68 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire67;
  reg signed [(4'hb):(1'h0)] reg66 = (1'h0);
  wire [(5'h13):(1'h0)] wire65;
  wire [(4'hb):(1'h0)] wire64;
  wire signed [(4'h8):(1'h0)] wire63;
  reg signed [(4'hc):(1'h0)] reg62 = (1'h0);
  reg [(5'h15):(1'h0)] reg61 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg60 = (1'h0);
  reg [(2'h2):(1'h0)] reg59 = (1'h0);
  reg [(4'hf):(1'h0)] reg58 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire57;
  reg [(4'hd):(1'h0)] reg56 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg55 = (1'h0);
  reg [(4'he):(1'h0)] reg54 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg53 = (1'h0);
  reg [(5'h10):(1'h0)] forvar52 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar51 = (1'h0);
  reg [(3'h5):(1'h0)] reg50 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire49;
  wire signed [(2'h3):(1'h0)] wire48;
  reg [(4'h9):(1'h0)] reg47 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg46 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg45 = (1'h0);
  reg [(3'h5):(1'h0)] forvar44 = (1'h0);
  reg [(3'h7):(1'h0)] reg43 = (1'h0);
  reg [(4'hb):(1'h0)] reg42 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg41 = (1'h0);
  reg [(5'h14):(1'h0)] reg40 = (1'h0);
  reg [(2'h3):(1'h0)] forvar39 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg38 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar33 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg37 = (1'h0);
  reg [(2'h3):(1'h0)] reg36 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg35 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg34 = (1'h0);
  reg [(4'hb):(1'h0)] reg33 = (1'h0);
  reg [(4'ha):(1'h0)] reg32 = (1'h0);
  reg [(5'h13):(1'h0)] reg31 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg30 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg29 = (1'h0);
  reg [(3'h6):(1'h0)] reg28 = (1'h0);
  reg [(5'h13):(1'h0)] reg27 = (1'h0);
  reg [(3'h7):(1'h0)] reg26 = (1'h0);
  reg [(4'he):(1'h0)] reg25 = (1'h0);
  reg [(3'h5):(1'h0)] reg24 = (1'h0);
  reg [(2'h3):(1'h0)] reg23 = (1'h0);
  reg [(4'hb):(1'h0)] reg22 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg21 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire20;
  reg [(5'h12):(1'h0)] reg19 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg18 = (1'h0);
  reg [(5'h15):(1'h0)] reg17 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg16 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg15 = (1'h0);
  reg [(4'he):(1'h0)] forvar14 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg13 = (1'h0);
  reg [(3'h7):(1'h0)] reg12 = (1'h0);
  reg [(4'h9):(1'h0)] reg11 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg10 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg9 = (1'h0);
  reg [(4'h9):(1'h0)] reg8 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar7 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5 = (1'h0);
  wire [(4'hb):(1'h0)] wire4;
  assign y = {wire461,
                 reg460,
                 reg459,
                 reg458,
                 forvar457,
                 reg456,
                 reg455,
                 forvar454,
                 reg453,
                 reg452,
                 wire450,
                 reg71,
                 reg70,
                 reg69,
                 forvar68,
                 wire67,
                 reg66,
                 wire65,
                 wire64,
                 wire63,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 wire57,
                 reg56,
                 reg55,
                 reg54,
                 reg53,
                 forvar52,
                 forvar51,
                 reg50,
                 wire49,
                 wire48,
                 reg47,
                 reg46,
                 reg45,
                 forvar44,
                 reg43,
                 reg42,
                 reg41,
                 reg40,
                 forvar39,
                 reg38,
                 forvar33,
                 reg37,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 reg32,
                 reg31,
                 reg30,
                 reg29,
                 reg28,
                 reg27,
                 reg26,
                 reg25,
                 reg24,
                 reg23,
                 reg22,
                 reg21,
                 wire20,
                 reg19,
                 reg18,
                 reg17,
                 reg16,
                 reg15,
                 forvar14,
                 reg13,
                 reg12,
                 reg11,
                 reg10,
                 reg9,
                 reg8,
                 forvar7,
                 reg6,
                 reg5,
                 wire4,
                 (1'h0)};
  assign wire4 = $unsigned(wire2[(4'hb):(3'h7)]);
  always
    @(posedge clk) begin
      reg5 <= {(^~$unsigned((~|(wire0 ? wire3 : wire1)))),
          $signed($signed(wire4[(3'h4):(1'h0)]))};
      reg6 <= $signed(wire1[(1'h0):(1'h0)]);
      for (forvar7 = (1'h0); (forvar7 < (2'h2)); forvar7 = (forvar7 + (1'h1)))
        begin
          reg8 <= (|($signed($unsigned((wire0 ? reg5 : (7'h42)))) ?
              wire1 : {$unsigned($signed(wire4))}));
          reg9 <= $unsigned(((8'h9f) <= wire3));
          reg10 <= {reg6, wire4};
          reg11 <= wire2;
        end
      reg12 <= ((reg9 + wire0[(3'h6):(2'h2)]) == $unsigned($signed(wire1[(3'h4):(3'h4)])));
    end
  always
    @(posedge clk) begin
      reg13 <= {reg12[(1'h1):(1'h0)],
          ((reg11[(1'h0):(1'h0)] ~^ (8'ha3)) ? reg8 : (8'ha6))};
      for (forvar14 = (1'h0); (forvar14 < (1'h0)); forvar14 = (forvar14 + (1'h1)))
        begin
          reg15 <= (((((reg11 ? forvar7 : forvar7) ~^ $unsigned(wire0)) ?
                  {forvar7[(1'h1):(1'h0)]} : $unsigned((~wire0))) ?
              $unsigned($unsigned((reg12 | reg9))) : reg8) * reg9);
          reg16 <= wire4;
        end
      reg17 = (reg15 ?
          ($unsigned(($unsigned(forvar7) > wire4[(2'h2):(1'h0)])) != (-(reg5[(4'ha):(3'h5)] - (wire2 ~^ (8'ha1))))) : $signed(reg12[(3'h4):(2'h3)]));
    end
  always
    @(posedge clk) begin
      reg18 <= $signed($unsigned($signed(reg16)));
      reg19 = (|({($signed((7'h42)) - {reg6, (8'h9c)}),
              (wire1 || $unsigned(reg10))} ?
          reg5 : (^~forvar7[(2'h2):(1'h0)])));
    end
  assign wire20 = reg18[(2'h2):(1'h0)];
  always
    @(posedge clk) begin
      reg21 <= wire20[(5'h11):(4'h9)];
      reg22 <= {{$unsigned($unsigned((wire1 ? reg9 : reg12))),
              $unsigned(((reg18 <<< forvar14) ? reg21 : $unsigned(reg17)))}};
      reg23 = (-$signed($unsigned((reg5 - (forvar14 ? reg22 : reg12)))));
      reg24 <= ($signed(reg12) ~^ (!($unsigned($signed(reg23)) * ({reg15,
              reg13} ?
          forvar14[(4'hb):(4'h8)] : (reg11 ? reg23 : wire2)))));
    end
  always
    @(posedge clk) begin
      reg25 <= (8'hb3);
      reg26 = (reg13[(4'h8):(3'h6)] < (^wire0[(3'h7):(3'h6)]));
      reg27 <= ($signed($signed((wire20 ? $unsigned(forvar7) : (^~reg11)))) ?
          (({$signed(reg25)} < ({reg13} <= reg26)) <= $signed((8'ha2))) : $unsigned((((~&wire1) ~^ wire1) >> $unsigned((reg18 ?
              reg26 : reg12)))));
      reg28 <= (8'ha9);
      reg29 <= reg27[(4'hd):(4'hd)];
    end
  always
    @(posedge clk) begin
      reg30 <= wire0;
      reg31 <= (&{reg6[(2'h2):(1'h0)], $signed(reg21[(3'h4):(2'h3)])});
      reg32 = ($unsigned((8'ha0)) ?
          $unsigned((7'h40)) : $unsigned($signed(wire3)));
      if (((($signed(reg32[(4'ha):(3'h7)]) < $signed((reg32 ?
              (8'ha2) : reg18))) - ($signed((reg22 * reg26)) >>> ($signed(reg18) < (wire0 <= wire20)))) ?
          (reg17[(5'h12):(4'hd)] ?
              forvar7[(1'h0):(1'h0)] : (+(!(+reg25)))) : {(|wire20),
              wire20[(3'h6):(1'h1)]}))
        begin
          reg33 <= (wire0 & $unsigned($signed((~|reg10[(3'h4):(3'h4)]))));
          reg34 = (reg13[(4'hd):(3'h4)] << (~|reg27));
          reg35 = (^reg24);
          reg36 <= (({(reg12 <= forvar7[(1'h1):(1'h1)]), {$unsigned((8'ha5))}} ?
              $unsigned(reg8) : ((+$unsigned(reg27)) ?
                  ((^reg18) << $unsigned((8'hba))) : (((7'h44) && reg19) ?
                      {(8'hb4)} : {reg29}))) - reg28[(2'h2):(1'h1)]);
          reg37 <= reg33[(1'h0):(1'h0)];
        end
      else
        begin
          for (forvar33 = (1'h0); (forvar33 < (2'h3)); forvar33 = (forvar33 + (1'h1)))
            begin
              reg34 <= (+{$signed((-(reg31 ^~ reg34)))});
              reg35 <= (wire2 ?
                  (!($signed((~^reg18)) ?
                      (8'ha3) : $signed((-reg10)))) : (~(8'ha2)));
              reg36 <= ($unsigned(wire1) ?
                  (~reg28[(2'h2):(1'h0)]) : {reg34[(4'h9):(4'h9)]});
              reg37 <= {reg10,
                  ($signed($signed((8'ha2))) ?
                      ($signed(reg6) ?
                          $signed({wire3}) : reg22) : (reg37[(2'h2):(1'h1)] & ((reg33 > reg10) | {reg31})))};
            end
          reg38 = reg30[(3'h4):(1'h1)];
        end
      for (forvar39 = (1'h0); (forvar39 < (1'h0)); forvar39 = (forvar39 + (1'h1)))
        begin
          reg40 = (reg28[(1'h1):(1'h0)] ?
              $signed((!({forvar33, reg33} ?
                  reg24[(3'h4):(3'h4)] : ((8'hac) << reg18)))) : (reg12[(1'h1):(1'h0)] ?
                  {$unsigned(forvar7)} : ((wire4[(4'ha):(4'ha)] == {(8'ha3)}) || $unsigned($signed(reg21)))));
          reg41 <= {(reg24 ?
                  $unsigned(forvar39) : (reg30[(3'h7):(1'h0)] >> (-reg33)))};
          reg42 = $unsigned(($signed((^reg12[(3'h6):(1'h1)])) != (^forvar33[(1'h1):(1'h0)])));
          reg43 <= $unsigned(reg23[(1'h0):(1'h0)]);
          for (forvar44 = (1'h0); (forvar44 < (2'h3)); forvar44 = (forvar44 + (1'h1)))
            begin
              reg45 <= $unsigned(({($signed(reg16) < (forvar7 ? reg11 : reg43)),
                  reg37} * ({(~reg24)} ?
                  $signed($signed(reg11)) : (~&{forvar14}))));
              reg46 <= $unsigned(reg32[(4'h9):(4'h8)]);
              reg47 = reg28[(3'h4):(3'h4)];
            end
        end
    end
  assign wire48 = (({reg30[(3'h6):(1'h0)]} ?
                      ({(reg31 ? reg36 : reg29)} ?
                          ($unsigned(reg38) == (^reg9)) : $unsigned(reg34)) : $signed((&$signed((8'hb2))))) ~^ $signed((-reg5)));
  assign wire49 = ($unsigned($unsigned((&(reg6 ?
                      reg37 : wire20)))) | ($unsigned((^$signed(reg22))) ?
                      reg8 : $unsigned((^(forvar7 ? reg32 : reg37)))));
  always
    @(posedge clk) begin
      reg50 <= $signed($signed({reg23[(2'h2):(1'h0)]}));
      for (forvar51 = (1'h0); (forvar51 < (2'h3)); forvar51 = (forvar51 + (1'h1)))
        begin
          for (forvar52 = (1'h0); (forvar52 < (1'h0)); forvar52 = (forvar52 + (1'h1)))
            begin
              reg53 <= $signed(wire3);
              reg54 <= $unsigned($signed((-(~&(reg9 == reg31)))));
            end
          reg55 <= $unsigned(reg36);
          reg56 <= reg36;
        end
    end
  assign wire57 = $signed($unsigned({wire4}));
  always
    @(posedge clk) begin
      reg58 = (+$signed(((wire0 ?
          $signed(reg56) : (!(8'had))) >>> $unsigned($unsigned(reg54)))));
      reg59 <= reg5[(2'h3):(1'h0)];
      reg60 = (wire49[(3'h6):(3'h4)] ?
          (($unsigned(reg30[(3'h4):(3'h4)]) + {reg47,
              (reg23 ?
                  reg35 : reg16)}) != $unsigned(((reg32 <<< reg42) * (8'ha7)))) : forvar52[(3'h6):(2'h2)]);
      reg61 <= (($unsigned(wire49[(2'h3):(2'h3)]) ?
              $unsigned($signed((wire49 ?
                  reg46 : reg35))) : ((|reg21) ~^ forvar52[(5'h10):(3'h4)])) ?
          reg26[(3'h5):(3'h4)] : $signed($signed(forvar51)));
      reg62 <= (((+(!reg58[(1'h1):(1'h1)])) >>> $signed(wire49)) & $signed((reg47[(3'h4):(3'h4)] != (+(wire4 ^~ reg29)))));
    end
  assign wire63 = reg60;
  assign wire64 = ({reg43} > {$signed($unsigned(reg24)), reg41[(4'hb):(2'h3)]});
  assign wire65 = (reg24[(3'h4):(1'h0)] >> ((reg17[(5'h13):(4'hc)] ?
                      $signed(reg28) : (wire64[(4'ha):(3'h5)] || reg27[(4'h9):(3'h7)])) || (reg42 ?
                      ($unsigned(reg23) ?
                          reg6[(4'h8):(1'h0)] : reg42) : $unsigned({reg9}))));
  always
    @(posedge clk) begin
      reg66 = (($unsigned($signed($signed(reg56))) ?
          forvar44 : ($signed($unsigned(reg46)) ?
              ((reg40 >= reg32) ?
                  reg34 : $signed((8'hab))) : reg43)) || (~|$signed($signed($unsigned((8'haa))))));
    end
  assign wire67 = (((((reg60 ?
                      wire64 : wire65) ^~ (8'hb2)) <= reg54[(4'ha):(3'h7)]) || (($signed(reg27) ?
                          {reg30} : $signed(reg18)) ?
                      (((8'h9d) >> reg13) ?
                          $unsigned(reg9) : reg45) : forvar39[(1'h1):(1'h0)])) * (8'h9f));
  always
    @(posedge clk) begin
      for (forvar68 = (1'h0); (forvar68 < (1'h0)); forvar68 = (forvar68 + (1'h1)))
        begin
          reg69 <= (~&($signed(wire4) ?
              forvar39 : $signed(((~&wire48) ^ wire63))));
        end
      reg70 <= reg28[(3'h6):(2'h2)];
      reg71 <= $signed((|(^~reg11)));
    end
  module72 modinst451 (.wire76(reg25), .y(wire450), .wire74(wire2), .wire75(wire1), .clk(clk), .wire73(reg30));
  always
    @(posedge clk) begin
      reg452 <= $unsigned($unsigned(wire65));
      reg453 = (reg34[(3'h6):(2'h3)] ~^ $unsigned($signed($unsigned((reg70 ?
          reg21 : wire3)))));
      for (forvar454 = (1'h0); (forvar454 < (2'h2)); forvar454 = (forvar454 + (1'h1)))
        begin
          reg455 <= reg453[(4'ha):(4'ha)];
          reg456 <= reg58[(3'h6):(1'h1)];
          for (forvar457 = (1'h0); (forvar457 < (1'h0)); forvar457 = (forvar457 + (1'h1)))
            begin
              reg458 = (-$unsigned(((~|reg47[(2'h3):(1'h0)]) << ((reg23 || reg11) ?
                  (reg47 <= reg13) : ((8'ha5) << reg26)))));
            end
        end
      reg459 <= reg69[(4'hb):(3'h7)];
      reg460 <= ($unsigned(($signed($unsigned(reg18)) ?
          reg24 : reg54[(2'h3):(2'h3)])) || reg23);
    end
  assign wire461 = $unsigned(reg12);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module72  (y, clk, wire73, wire74, wire75, wire76);
  output wire [(32'h35c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire73;
  input wire signed [(4'hf):(1'h0)] wire74;
  input wire [(4'h8):(1'h0)] wire75;
  input wire [(4'he):(1'h0)] wire76;
  reg signed [(5'h14):(1'h0)] reg77 = (1'h0);
  reg [(5'h14):(1'h0)] reg78 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg79 = (1'h0);
  reg [(3'h6):(1'h0)] forvar80 = (1'h0);
  reg [(2'h2):(1'h0)] reg81 = (1'h0);
  reg [(4'hf):(1'h0)] reg82 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar83 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg84 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg85 = (1'h0);
  reg [(5'h14):(1'h0)] reg86 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg87 = (1'h0);
  reg [(4'hb):(1'h0)] reg88 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar89 = (1'h0);
  reg signed [(4'he):(1'h0)] reg90 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar91 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg92 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg93 = (1'h0);
  reg [(4'h9):(1'h0)] reg94 = (1'h0);
  reg [(5'h15):(1'h0)] reg95 = (1'h0);
  reg [(4'hb):(1'h0)] reg96 = (1'h0);
  reg [(3'h7):(1'h0)] reg97 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg98 = (1'h0);
  reg [(5'h14):(1'h0)] reg99 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg100 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg101 = (1'h0);
  reg [(2'h3):(1'h0)] forvar102 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg103 = (1'h0);
  reg [(4'ha):(1'h0)] reg104 = (1'h0);
  reg signed [(4'he):(1'h0)] reg105 = (1'h0);
  reg [(5'h12):(1'h0)] forvar106 = (1'h0);
  reg [(5'h11):(1'h0)] reg107 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg108 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg109 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg110 = (1'h0);
  reg [(5'h10):(1'h0)] reg111 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg112 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg113 = (1'h0);
  reg [(3'h7):(1'h0)] reg114 = (1'h0);
  reg [(5'h10):(1'h0)] reg115 = (1'h0);
  reg [(4'hb):(1'h0)] reg116 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire117;
  reg signed [(3'h4):(1'h0)] forvar118 = (1'h0);
  reg [(5'h10):(1'h0)] reg119 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg120 = (1'h0);
  reg [(5'h13):(1'h0)] reg121 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg122 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg123 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg124 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg125 = (1'h0);
  reg [(4'ha):(1'h0)] reg126 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg127 = (1'h0);
  reg [(3'h7):(1'h0)] reg128 = (1'h0);
  wire [(3'h6):(1'h0)] wire129;
  wire signed [(4'h8):(1'h0)] wire130;
  wire [(3'h7):(1'h0)] wire207;
  wire [(5'h15):(1'h0)] wire209;
  wire [(5'h15):(1'h0)] wire210;
  reg signed [(5'h10):(1'h0)] forvar211 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg212 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg213 = (1'h0);
  reg [(5'h15):(1'h0)] reg214 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg215 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar216 = (1'h0);
  reg [(5'h12):(1'h0)] reg217 = (1'h0);
  reg [(5'h12):(1'h0)] reg218 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg219 = (1'h0);
  reg [(4'hc):(1'h0)] reg220 = (1'h0);
  reg [(4'hc):(1'h0)] reg221 = (1'h0);
  wire [(5'h15):(1'h0)] wire448;
  assign y = {reg77,
                 reg78,
                 reg79,
                 forvar80,
                 reg81,
                 reg82,
                 forvar83,
                 reg84,
                 reg85,
                 reg86,
                 reg87,
                 reg88,
                 forvar89,
                 reg90,
                 forvar91,
                 reg92,
                 reg93,
                 reg94,
                 reg95,
                 reg96,
                 reg97,
                 reg98,
                 reg99,
                 reg100,
                 reg101,
                 forvar102,
                 reg103,
                 reg104,
                 reg105,
                 forvar106,
                 reg107,
                 reg108,
                 reg109,
                 reg110,
                 reg111,
                 reg112,
                 reg113,
                 reg114,
                 reg115,
                 reg116,
                 wire117,
                 forvar118,
                 reg119,
                 reg120,
                 reg121,
                 reg122,
                 reg123,
                 reg124,
                 reg125,
                 reg126,
                 reg127,
                 reg128,
                 wire129,
                 wire130,
                 wire207,
                 wire209,
                 wire210,
                 forvar211,
                 reg212,
                 reg213,
                 reg214,
                 reg215,
                 forvar216,
                 reg217,
                 reg218,
                 reg219,
                 reg220,
                 reg221,
                 wire448,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg77 = wire75[(3'h4):(2'h3)];
      reg78 <= (wire76 ? $signed($signed((~&(wire74 ~^ wire76)))) : wire76);
      reg79 <= ((^$signed($unsigned(wire75[(3'h5):(1'h0)]))) ?
          $signed($unsigned((wire74 ? wire76 : $unsigned(wire73)))) : reg78);
    end
  always
    @(posedge clk) begin
      for (forvar80 = (1'h0); (forvar80 < (2'h3)); forvar80 = (forvar80 + (1'h1)))
        begin
          reg81 = $signed({(((reg77 ? forvar80 : wire76) ?
                  $signed(wire73) : $signed(wire75)) > (8'ha9))});
          reg82 <= reg81[(2'h2):(2'h2)];
          for (forvar83 = (1'h0); (forvar83 < (3'h4)); forvar83 = (forvar83 + (1'h1)))
            begin
              reg84 <= wire75[(2'h3):(2'h3)];
              reg85 <= ((((~|(reg82 ? wire76 : reg84)) <<< ((forvar80 ?
                          forvar80 : wire73) ?
                      (forvar80 ? (7'h44) : reg84) : (-(7'h41)))) ?
                  $signed($signed((&wire75))) : ((forvar83[(3'h5):(2'h3)] ?
                          $signed(reg77) : (forvar83 != reg84)) ?
                      (8'hb0) : wire73)) >= $signed($signed((~^$unsigned(reg82)))));
              reg86 <= $unsigned((^$unsigned($unsigned($signed(reg81)))));
            end
          reg87 <= wire73;
          reg88 = (($unsigned(wire73) ?
              ($unsigned((reg85 * (8'hb1))) ?
                  (forvar83[(1'h0):(1'h0)] | (^reg77)) : reg85) : $signed((wire73[(3'h6):(3'h5)] ?
                  (8'ha6) : ((7'h43) & reg81)))) >= reg87[(2'h2):(2'h2)]);
        end
      for (forvar89 = (1'h0); (forvar89 < (2'h2)); forvar89 = (forvar89 + (1'h1)))
        begin
          reg90 = $signed((reg88 ?
              $unsigned((((8'hb5) >> reg81) >> (wire76 ?
                  forvar80 : reg85))) : forvar89[(3'h4):(3'h4)]));
          for (forvar91 = (1'h0); (forvar91 < (3'h4)); forvar91 = (forvar91 + (1'h1)))
            begin
              reg92 <= ($signed(forvar83) * (^wire76));
            end
          if (wire75[(3'h4):(2'h3)])
            begin
              reg93 = reg87;
              reg94 = $unsigned(reg90[(3'h5):(3'h5)]);
              reg95 <= $unsigned(wire76);
            end
          else
            begin
              reg93 <= reg82;
              reg94 = $unsigned($unsigned($unsigned($signed(reg93))));
              reg95 = (&$signed(($signed((reg87 ?
                  (8'ha3) : wire75)) > $signed(reg87[(2'h3):(1'h1)]))));
              reg96 <= ((^~forvar80[(3'h6):(3'h6)]) ~^ $unsigned($signed($unsigned(forvar83))));
            end
          reg97 = reg86;
          reg98 <= (reg93 ~^ (^($signed($signed(wire73)) ?
              ($signed(reg95) < $signed(reg96)) : $signed($unsigned(forvar83)))));
        end
    end
  always
    @(posedge clk) begin
      reg99 <= ((reg77[(4'h9):(2'h3)] > $unsigned(($signed((8'ha7)) == (^~reg96)))) ?
          $unsigned($unsigned(($signed(reg87) ?
              $unsigned(reg95) : (wire73 ? reg85 : reg87)))) : (^reg78));
      reg100 <= $signed($signed($signed({$unsigned(wire75)})));
      reg101 <= ($unsigned(((^~wire73) >>> $signed({reg90, reg98}))) ?
          (~^((wire75[(1'h1):(1'h1)] ?
              (~reg95) : reg99) != $signed((reg88 & reg88)))) : {($unsigned($unsigned(reg95)) ?
                  reg95 : reg97[(3'h4):(3'h4)])});
      for (forvar102 = (1'h0); (forvar102 < (2'h2)); forvar102 = (forvar102 + (1'h1)))
        begin
          reg103 = reg84[(2'h3):(2'h3)];
          reg104 = $signed((^~$signed($signed((&(8'ha2))))));
          reg105 <= $signed((~|reg84[(2'h2):(1'h1)]));
          for (forvar106 = (1'h0); (forvar106 < (1'h0)); forvar106 = (forvar106 + (1'h1)))
            begin
              reg107 <= reg105;
            end
          reg108 <= (~|((((wire73 ^~ forvar102) == (forvar91 <<< forvar102)) ?
                  $unsigned({reg90, forvar83}) : {((8'h9c) ?
                          (8'ha5) : wire75)}) ?
              $unsigned($signed((wire73 ?
                  reg97 : reg82))) : $unsigned({(~(8'hb8))})));
        end
      reg109 <= wire73;
    end
  always
    @(posedge clk) begin
      reg110 <= ((reg107 ?
          $unsigned($unsigned(reg100[(3'h4):(1'h0)])) : (reg96 - (wire74[(4'hf):(1'h1)] ?
              (~^reg87) : reg86))) == (8'hb6));
      reg111 <= reg90;
      reg112 <= {($unsigned((8'hae)) ?
              (reg79[(3'h4):(3'h4)] && (reg94[(2'h2):(1'h1)] ?
                  (+reg85) : (!(8'ha7)))) : $signed($unsigned(reg94)))};
      reg113 <= (8'h9d);
    end
  always
    @(posedge clk) begin
      reg114 <= (wire73 ^~ (!reg112[(3'h7):(3'h5)]));
    end
  always
    @(posedge clk) begin
      reg115 <= (wire76 ? (8'hb3) : (-$signed(reg100)));
    end
  always
    @(posedge clk) begin
      reg116 <= ($unsigned({(~&reg84[(1'h1):(1'h0)]),
          (wire73 ?
              $signed(reg100) : $unsigned(reg101))}) <<< {$unsigned($signed($unsigned(reg90))),
          (~&$signed(((7'h40) << reg104)))});
    end
  assign wire117 = ((($signed(wire75) ?
                       ((reg92 ?
                           reg90 : forvar91) <<< (~|reg101)) : (~&$unsigned(reg101))) * {((^reg86) ?
                           (reg88 < reg88) : $signed(reg110)),
                       $signed({(8'haa)})}) >>> $signed((~(8'ha4))));
  always
    @(posedge clk) begin
      for (forvar118 = (1'h0); (forvar118 < (2'h3)); forvar118 = (forvar118 + (1'h1)))
        begin
          reg119 = (-reg81[(1'h0):(1'h0)]);
          reg120 <= $unsigned($signed($unsigned(($unsigned(reg84) ?
              $unsigned(reg86) : (reg79 > forvar89)))));
          reg121 = ($signed((^~(^~$signed(reg86)))) && $signed(reg86));
        end
      reg122 <= ((^$signed(reg81[(1'h1):(1'h0)])) ^ ($unsigned(($unsigned(reg81) ^ (wire73 ?
              reg81 : reg107))) ?
          $unsigned(reg95[(4'hf):(4'hb)]) : wire76));
      reg123 = {reg84, $unsigned($unsigned({(forvar118 >> reg103)}))};
      reg124 <= reg79[(3'h5):(3'h4)];
    end
  always
    @(posedge clk) begin
      reg125 <= $unsigned($unsigned((((reg88 & reg77) ?
              $signed((8'hba)) : reg109) ?
          ($unsigned(reg100) ?
              reg94[(2'h2):(1'h1)] : (^~reg111)) : (reg108 ^ (|forvar91)))));
      reg126 <= (reg105 ?
          forvar118 : $unsigned({$unsigned((forvar89 ^~ (8'ha2))),
              ($signed(reg114) >> reg107)}));
      reg127 <= ($unsigned((reg82 + (((8'ha6) ? reg121 : forvar89) ?
          reg104 : (8'ha8)))) >> $unsigned($unsigned({$unsigned(reg105)})));
    end
  always
    @(posedge clk) begin
      reg128 = $unsigned(reg78);
    end
  assign wire129 = ($unsigned($unsigned(reg90[(2'h3):(1'h1)])) ?
                       (reg125 ?
                           ((&(~^reg97)) ?
                               (!(&reg103)) : (reg98 | $unsigned(reg84))) : reg100) : (-reg92[(4'hb):(3'h6)]));
  assign wire130 = (&($unsigned((~^reg87)) ?
                       $signed((^~(reg114 ?
                           (8'ha5) : reg98))) : (^($unsigned(reg87) ?
                           ((8'hab) ?
                               forvar89 : (8'hb8)) : reg128[(1'h0):(1'h0)]))));
  module131 modinst208 (wire207, clk, reg86, reg119, reg92, reg107);
  assign wire209 = $signed((reg110 ?
                       {((reg81 && (8'ha9)) & (wire76 ? reg123 : forvar89)),
                           (reg123[(3'h4):(3'h4)] ?
                               forvar89[(3'h4):(3'h4)] : (reg116 == reg98))} : forvar102));
  assign wire210 = ($unsigned(reg94[(3'h7):(3'h7)]) ?
                       $unsigned((reg95[(3'h5):(3'h5)] ?
                           ($unsigned(reg125) ?
                               ((8'h9f) ?
                                   reg125 : wire74) : reg85[(4'hd):(4'h9)]) : ((8'hbf) >> $signed((7'h40))))) : $unsigned({((~^reg87) >>> $signed(forvar80)),
                           $signed((forvar118 ? forvar106 : forvar118))}));
  always
    @(posedge clk) begin
      for (forvar211 = (1'h0); (forvar211 < (3'h4)); forvar211 = (forvar211 + (1'h1)))
        begin
          reg212 <= (wire209[(4'hf):(1'h0)] || $unsigned((((~|reg127) ?
                  $unsigned(forvar118) : (-reg126)) ?
              reg108 : (&$unsigned(reg113)))));
          reg213 <= (~|$unsigned({reg100[(1'h0):(1'h0)]}));
          reg214 <= $signed(reg97[(3'h7):(1'h0)]);
          reg215 <= ($signed($signed(reg126)) ^~ (((wire73[(1'h0):(1'h0)] << $signed(reg86)) >>> reg126[(1'h0):(1'h0)]) ?
              reg120 : $signed(($signed(reg213) ?
                  {forvar91, wire76} : (^reg119)))));
          for (forvar216 = (1'h0); (forvar216 < (1'h1)); forvar216 = (forvar216 + (1'h1)))
            begin
              reg217 <= (wire74 ?
                  ((8'h9f) ? reg96[(3'h4):(1'h1)] : reg112) : wire74);
              reg218 <= reg109[(3'h5):(3'h5)];
            end
        end
      reg219 = ($unsigned($signed($signed($unsigned(wire210)))) ^~ $unsigned(((reg217[(5'h10):(3'h5)] ?
          reg81 : $unsigned(forvar118)) * $unsigned((&reg215)))));
      reg220 <= wire130[(2'h2):(1'h1)];
      reg221 <= $unsigned((reg103 & $unsigned($unsigned(((8'hbf) ?
          wire76 : (7'h41))))));
    end
  module222 modinst449 (.wire225(forvar89), .wire226(reg78), .y(wire448), .wire224(wire210), .wire223(reg82), .clk(clk), .wire227(reg96));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module222
#( parameter param446 = (({(^~{(8'ha4)})} ? (~|{((8'hb4) << (8'hb3)), (|(7'h40))}) : (&((8'hae) >= ((7'h41) ? (8'hbe) : (8'hab))))) ? ((~&(~(~^(8'ha6)))) | (((-(8'haf)) <<< (^(8'ha5))) ? (((7'h41) ? (8'hb4) : (8'hb3)) ? (&(8'h9d)) : (+(8'ha5))) : ({(8'hab), (8'had)} == ((8'hbb) ? (8'hb1) : (8'hb0))))) : (((|((8'hac) + (8'ha5))) == (+(~&(8'ha7)))) ? ({(~^(8'h9c)), ((8'haf) ? (8'hab) : (7'h44))} ? {{(8'hb8)}, ((8'ha5) ? (7'h41) : (8'hbf))} : (((8'ha2) ^~ (8'hb0)) || (8'ha6))) : ((((7'h42) <<< (8'hb3)) ^~ ((8'hb4) ? (8'ha3) : (8'hba))) | ({(8'haa), (8'hb3)} ? (-(8'hbb)) : ((8'hab) & (8'hbf))))))
, parameter param447 = (({(param446 >= (~param446))} ? param446 : param446) ? (param446 > param446) : {param446}) )
(y, clk, wire223, wire224, wire225, wire226, wire227);
  output wire [(32'h1d3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire223;
  input wire signed [(5'h15):(1'h0)] wire224;
  input wire signed [(4'hc):(1'h0)] wire225;
  input wire [(5'h14):(1'h0)] wire226;
  input wire [(4'hb):(1'h0)] wire227;
  wire [(4'hc):(1'h0)] wire445;
  wire signed [(4'h9):(1'h0)] wire444;
  reg [(4'h9):(1'h0)] reg443 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg442 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg441 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg440 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg228 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg229 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg230 = (1'h0);
  reg [(3'h5):(1'h0)] reg231 = (1'h0);
  reg [(5'h11):(1'h0)] forvar232 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg233 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar234 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg235 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg236 = (1'h0);
  reg [(4'h9):(1'h0)] reg237 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg238 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar239 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg240 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg241 = (1'h0);
  reg signed [(4'he):(1'h0)] reg242 = (1'h0);
  reg [(4'he):(1'h0)] reg243 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg244 = (1'h0);
  reg [(3'h4):(1'h0)] reg245 = (1'h0);
  wire [(2'h3):(1'h0)] wire246;
  reg signed [(3'h6):(1'h0)] reg247 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg248 = (1'h0);
  reg [(5'h10):(1'h0)] forvar249 = (1'h0);
  reg [(3'h4):(1'h0)] reg250 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg251 = (1'h0);
  reg [(4'he):(1'h0)] reg252 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire253;
  wire [(4'h9):(1'h0)] wire419;
  wire signed [(5'h14):(1'h0)] wire421;
  wire signed [(4'h9):(1'h0)] wire422;
  reg [(2'h3):(1'h0)] reg423 = (1'h0);
  reg [(4'h9):(1'h0)] reg424 = (1'h0);
  wire [(5'h13):(1'h0)] wire425;
  wire signed [(3'h5):(1'h0)] wire426;
  wire [(2'h3):(1'h0)] wire438;
  assign y = {wire445,
                 wire444,
                 reg443,
                 reg442,
                 reg441,
                 reg440,
                 reg228,
                 reg229,
                 reg230,
                 reg231,
                 forvar232,
                 reg233,
                 forvar234,
                 reg235,
                 reg236,
                 reg237,
                 reg238,
                 forvar239,
                 reg240,
                 reg241,
                 reg242,
                 reg243,
                 reg244,
                 reg245,
                 wire246,
                 reg247,
                 reg248,
                 forvar249,
                 reg250,
                 reg251,
                 reg252,
                 wire253,
                 wire419,
                 wire421,
                 wire422,
                 reg423,
                 reg424,
                 wire425,
                 wire426,
                 wire438,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg228 <= $unsigned(wire223);
      reg229 = $signed($unsigned($unsigned({(^wire224), $unsigned(wire224)})));
    end
  always
    @(posedge clk) begin
      reg230 <= $unsigned($unsigned(reg229[(4'h9):(3'h5)]));
      reg231 <= {((~wire226) ?
              {wire226[(4'ha):(3'h4)]} : (^~((~^(8'had)) <<< wire226)))};
      for (forvar232 = (1'h0); (forvar232 < (1'h0)); forvar232 = (forvar232 + (1'h1)))
        begin
          reg233 <= reg231;
          for (forvar234 = (1'h0); (forvar234 < (3'h4)); forvar234 = (forvar234 + (1'h1)))
            begin
              reg235 <= reg229[(2'h2):(2'h2)];
              reg236 <= reg229;
              reg237 <= $unsigned(wire225[(4'hb):(3'h4)]);
              reg238 <= $signed((^(~&reg236[(3'h4):(2'h2)])));
            end
          for (forvar239 = (1'h0); (forvar239 < (3'h4)); forvar239 = (forvar239 + (1'h1)))
            begin
              reg240 <= (reg233[(3'h6):(2'h2)] ?
                  ({(8'hb0)} | $signed((~|wire225))) : reg233);
              reg241 <= wire226[(4'h8):(1'h1)];
              reg242 = wire225[(2'h3):(2'h3)];
              reg243 = ($signed(wire227[(3'h5):(1'h0)]) ?
                  wire226[(1'h0):(1'h0)] : $signed(((8'hbe) ?
                      reg233 : ($signed(wire224) ?
                          reg241[(1'h1):(1'h1)] : (reg241 ?
                              reg240 : (8'ha9))))));
              reg244 = ($signed($unsigned((wire227 ?
                      {reg236} : (reg233 || wire227)))) ?
                  (wire224 ?
                      (&wire224[(5'h11):(4'hf)]) : (wire223[(4'hb):(3'h4)] ?
                          {(~wire223)} : (|(forvar239 ?
                              reg243 : reg240)))) : (forvar232[(5'h10):(4'he)] + $unsigned(forvar232)));
            end
          reg245 <= wire227;
        end
    end
  assign wire246 = $signed((($unsigned(((8'hac) ?
                       reg233 : wire227)) ^ (reg242[(4'hb):(3'h5)] ?
                       $unsigned(reg240) : (8'hab))) <= wire225[(4'hc):(4'ha)]));
  always
    @(posedge clk) begin
      reg247 <= $signed(wire227[(4'hb):(1'h1)]);
      reg248 <= $signed((wire227[(1'h0):(1'h0)] ?
          ((~^reg240[(3'h4):(3'h4)]) != (!reg235[(3'h5):(1'h1)])) : $unsigned((forvar232 ?
              (8'ha9) : $signed(wire223)))));
      for (forvar249 = (1'h0); (forvar249 < (1'h0)); forvar249 = (forvar249 + (1'h1)))
        begin
          reg250 = $signed((reg237 != $unsigned(((reg241 | forvar249) ?
              {reg247, reg237} : (-reg229)))));
        end
      reg251 <= {reg241};
      reg252 <= (wire246 ^~ (&{$signed((|(8'ha0))), {reg233[(1'h0):(1'h0)]}}));
    end
  assign wire253 = ($signed((((|(8'had)) <<< $unsigned(reg252)) ^ wire246[(1'h1):(1'h0)])) & ((8'had) ?
                       {$signed(reg235[(1'h1):(1'h0)])} : $unsigned(reg244)));
  module254 modinst420 (.wire257(forvar232), .y(wire419), .wire255(reg248), .wire258(reg235), .clk(clk), .wire256(reg244));
  assign wire421 = (~$unsigned(($unsigned(reg231) * (^$unsigned(reg243)))));
  assign wire422 = $unsigned($unsigned(reg233));
  always
    @(posedge clk) begin
      reg423 <= ((|(+reg238[(4'h8):(3'h6)])) ?
          (7'h41) : $signed($unsigned(($signed(reg230) ^~ (~&reg251)))));
      reg424 <= (({forvar232[(4'hc):(1'h1)]} + $signed(reg233[(4'h8):(3'h5)])) ?
          $unsigned({($signed(reg247) ? $signed(reg235) : (reg236 <<< wire253)),
              ($unsigned(wire421) > (reg240 + reg242))}) : ($signed(((!reg245) ^ (wire422 ~^ (7'h42)))) ?
              ($unsigned($unsigned(reg236)) || reg245) : ($signed(wire224[(5'h15):(2'h2)]) ?
                  $signed((wire224 >> wire422)) : $unsigned($unsigned(wire246)))));
    end
  assign wire425 = (wire246[(1'h0):(1'h0)] + $signed($unsigned({(|(8'ha0))})));
  assign wire426 = $signed((!$signed(reg240)));
  module427 modinst439 (wire438, clk, wire421, reg233, wire227, wire224, reg240);
  always
    @(posedge clk) begin
      reg440 = (($signed((reg244[(1'h0):(1'h0)] >= wire224)) ?
              $signed((reg248[(4'h8):(3'h6)] ~^ reg242[(2'h2):(2'h2)])) : reg244[(2'h2):(1'h0)]) ?
          wire227 : (|(^~$unsigned(reg240))));
      reg441 <= $signed(reg248);
    end
  always
    @(posedge clk) begin
      reg442 <= (((&$signed((-reg228))) ?
              {((~&reg231) ? {reg238, reg242} : (reg244 ? (8'haa) : (8'hac))),
                  (reg424 + (reg423 < (8'hb1)))} : (~&$unsigned(((8'ha6) ?
                  reg228 : reg228)))) ?
          (!wire227[(3'h7):(3'h5)]) : ($signed((-(reg248 ?
              forvar239 : forvar232))) ^~ forvar239));
      reg443 <= {(reg229[(4'h9):(4'h9)] ?
              (^wire421) : $signed($signed((!reg229)))),
          ({reg242[(4'h8):(3'h6)]} ?
              (((wire227 + (7'h44)) <= (~|reg440)) && reg235) : (reg248[(2'h2):(2'h2)] ^ wire224[(5'h10):(4'hb)]))};
    end
  assign wire444 = $unsigned($signed(wire425));
  assign wire445 = reg244;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module131  (y, clk, wire135, wire134, wire133, wire132);
  output wire [(32'ha5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire135;
  input wire signed [(5'h10):(1'h0)] wire134;
  input wire signed [(5'h15):(1'h0)] wire133;
  input wire signed [(5'h11):(1'h0)] wire132;
  reg [(4'he):(1'h0)] reg206 = (1'h0);
  reg [(3'h7):(1'h0)] reg205 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg204 = (1'h0);
  reg [(5'h10):(1'h0)] reg203 = (1'h0);
  wire [(5'h12):(1'h0)] wire202;
  wire signed [(5'h12):(1'h0)] wire201;
  reg signed [(4'hb):(1'h0)] reg200 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg199 = (1'h0);
  reg signed [(4'he):(1'h0)] reg198 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire196;
  wire signed [(4'h8):(1'h0)] wire159;
  wire [(2'h3):(1'h0)] wire158;
  wire [(4'h9):(1'h0)] wire157;
  wire signed [(5'h13):(1'h0)] wire155;
  assign y = {reg206,
                 reg205,
                 reg204,
                 reg203,
                 wire202,
                 wire201,
                 reg200,
                 reg199,
                 reg198,
                 wire196,
                 wire159,
                 wire158,
                 wire157,
                 wire155,
                 (1'h0)};
  module136 modinst156 (.wire139(wire135), .wire137(wire132), .wire140(wire133), .y(wire155), .clk(clk), .wire138(wire134));
  assign wire157 = (wire135 + wire132[(4'h8):(3'h5)]);
  assign wire158 = (7'h43);
  assign wire159 = ((~^$signed(($signed((8'hab)) ?
                       (wire157 << (8'ha8)) : wire158))) == ($signed(wire132[(5'h11):(4'hb)]) != wire157));
  module160 modinst197 (.wire162(wire132), .y(wire196), .wire164(wire134), .clk(clk), .wire161(wire135), .wire163(wire155));
  always
    @(posedge clk) begin
      reg198 = $unsigned({$unsigned(wire135),
          (wire196 >>> $unsigned((wire157 || wire159)))});
      reg199 = ((~&$unsigned({$unsigned(wire155)})) && (((wire134[(4'he):(3'h7)] == {wire132}) != ($unsigned(wire134) < $signed(wire133))) ^~ (^~(wire155[(1'h0):(1'h0)] <= (wire157 == wire155)))));
      reg200 <= (reg199[(4'hb):(3'h4)] ?
          (wire155[(3'h6):(3'h5)] ?
              wire157 : (wire132 ? (8'hab) : (&$signed((7'h44))))) : wire157);
    end
  assign wire201 = {((wire134 | $signed($signed(reg198))) >> $unsigned((8'ha0)))};
  assign wire202 = $signed($unsigned(({$unsigned(reg199)} - $signed(reg199[(2'h3):(2'h2)]))));
  always
    @(posedge clk) begin
      reg203 <= ($unsigned(wire155) ?
          ((|({wire134} * (wire133 ?
              reg198 : wire155))) >= $signed(wire158[(1'h0):(1'h0)])) : $unsigned($signed($unsigned((8'hb0)))));
      reg204 <= wire202;
      reg205 <= $unsigned($signed($signed((-(wire159 ? reg200 : reg200)))));
    end
  always
    @(posedge clk) begin
      reg206 <= $signed($signed((&$unsigned((~^reg205)))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module160
#( parameter param194 = ((+((8'ha2) ? ({(8'hab)} == (~^(8'ha7))) : (((8'h9e) <<< (8'ha7)) << ((8'hb3) <= (8'ha3))))) ? ({(^~{(8'hac), (8'hb8)})} <<< (({(8'hac)} ? (8'ha1) : ((7'h44) ? (8'hbd) : (8'ha9))) != (((7'h40) & (8'ha1)) ~^ ((8'ha0) ? (8'ha8) : (8'ha3))))) : (({{(8'ha2)}, ((8'hbb) ? (8'haf) : (8'hae))} >> (&((8'h9d) ? (8'hba) : (8'hb0)))) ^ ({(~|(8'hbb)), (!(8'hab))} ? ({(8'hb1)} ? ((8'ha0) ? (8'haa) : (8'hab)) : {(8'hac), (8'hb4)}) : {{(7'h41)}})))
, parameter param195 = param194 )
(y, clk, wire164, wire163, wire162, wire161);
  output wire [(32'h17a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire164;
  input wire [(5'h13):(1'h0)] wire163;
  input wire [(4'hc):(1'h0)] wire162;
  input wire [(5'h14):(1'h0)] wire161;
  wire signed [(4'he):(1'h0)] wire193;
  reg [(4'hf):(1'h0)] reg189 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar186 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg185 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg192 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg191 = (1'h0);
  reg [(5'h14):(1'h0)] reg190 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar189 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg188 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg187 = (1'h0);
  reg [(2'h3):(1'h0)] reg186 = (1'h0);
  reg [(4'h8):(1'h0)] forvar185 = (1'h0);
  reg [(4'hf):(1'h0)] reg184 = (1'h0);
  reg [(5'h10):(1'h0)] reg183 = (1'h0);
  reg [(5'h10):(1'h0)] reg182 = (1'h0);
  reg [(4'ha):(1'h0)] reg181 = (1'h0);
  reg [(5'h15):(1'h0)] forvar180 = (1'h0);
  reg signed [(4'he):(1'h0)] reg179 = (1'h0);
  reg [(2'h3):(1'h0)] reg178 = (1'h0);
  reg [(4'hb):(1'h0)] reg177 = (1'h0);
  reg [(3'h4):(1'h0)] reg176 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg175 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg174 = (1'h0);
  reg [(5'h11):(1'h0)] forvar173 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg172 = (1'h0);
  reg [(3'h6):(1'h0)] reg171 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar170 = (1'h0);
  reg [(4'hc):(1'h0)] reg169 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire168;
  wire signed [(4'h8):(1'h0)] wire167;
  wire [(4'hd):(1'h0)] wire166;
  wire signed [(5'h15):(1'h0)] wire165;
  assign y = {wire193,
                 reg189,
                 forvar186,
                 reg185,
                 reg192,
                 reg191,
                 reg190,
                 forvar189,
                 reg188,
                 reg187,
                 reg186,
                 forvar185,
                 reg184,
                 reg183,
                 reg182,
                 reg181,
                 forvar180,
                 reg179,
                 reg178,
                 reg177,
                 reg176,
                 reg175,
                 reg174,
                 forvar173,
                 reg172,
                 reg171,
                 forvar170,
                 reg169,
                 wire168,
                 wire167,
                 wire166,
                 wire165,
                 (1'h0)};
  assign wire165 = ($unsigned($signed($signed(wire163))) ~^ wire163);
  assign wire166 = $signed(((((wire164 >> wire164) | wire165) ?
                           (&wire163[(3'h4):(2'h3)]) : ((wire165 >> wire162) ^~ $signed(wire165))) ?
                       wire164[(1'h1):(1'h0)] : wire164));
  assign wire167 = $signed((wire161[(4'hd):(4'hb)] > (((wire163 ?
                           wire162 : (8'haf)) > (wire164 ^~ wire166)) ?
                       (wire165[(3'h6):(3'h5)] ?
                           (wire165 << wire166) : wire164) : $signed($unsigned(wire161)))));
  assign wire168 = wire161[(5'h11):(3'h7)];
  always
    @(posedge clk) begin
      reg169 <= $unsigned(wire166);
      for (forvar170 = (1'h0); (forvar170 < (1'h0)); forvar170 = (forvar170 + (1'h1)))
        begin
          reg171 <= wire162[(2'h2):(1'h1)];
          reg172 <= $unsigned($unsigned((wire161 >> $signed((!wire163)))));
          for (forvar173 = (1'h0); (forvar173 < (1'h1)); forvar173 = (forvar173 + (1'h1)))
            begin
              reg174 = (~|$signed((~$signed($unsigned((8'hb6))))));
              reg175 <= (($unsigned(wire166[(1'h1):(1'h1)]) ~^ ((8'h9f) ?
                      ($signed(wire166) ?
                          reg171 : $unsigned(reg174)) : $unsigned(wire161[(5'h10):(3'h6)]))) ?
                  ((reg174 ^~ wire162) || (~wire165[(5'h10):(4'hc)])) : wire162);
              reg176 <= ($unsigned((8'had)) ?
                  wire164[(5'h10):(4'hb)] : wire164[(4'hf):(4'h9)]);
              reg177 = (+($signed($unsigned((reg174 ? wire161 : forvar173))) ?
                  ($signed((|forvar173)) || $signed((~^wire168))) : wire164));
            end
          reg178 <= wire167;
        end
      reg179 <= ($signed(forvar170[(3'h6):(3'h6)]) <= ($unsigned($unsigned(reg171[(3'h6):(3'h4)])) ?
          ($signed($unsigned(reg178)) ?
              reg171 : reg175) : ($unsigned($signed(reg169)) ^ ((reg178 && wire166) + wire162[(3'h7):(2'h2)]))));
      for (forvar180 = (1'h0); (forvar180 < (2'h3)); forvar180 = (forvar180 + (1'h1)))
        begin
          if ((^(~^$unsigned((wire167 ? {forvar170, (8'ha5)} : wire162)))))
            begin
              reg181 <= (~^{wire161});
              reg182 <= $signed(($signed($unsigned({reg178,
                  wire168})) && (reg178[(2'h2):(1'h1)] & reg178)));
            end
          else
            begin
              reg181 <= ($unsigned(wire168) ?
                  $unsigned({((reg171 ? (8'hb1) : wire165) ?
                          {reg176} : reg176[(1'h1):(1'h0)])}) : (($signed((reg171 - (7'h40))) ?
                      (~(^forvar170)) : (^~$signed(wire166))) - (|reg176[(1'h1):(1'h1)])));
              reg182 <= {{(wire165 ?
                          {$unsigned(reg182),
                              $signed((8'hb7))} : ((forvar180 ^~ wire162) ?
                              $unsigned((8'hb7)) : (~^reg179))),
                      (!($signed(reg171) ?
                          reg176[(1'h1):(1'h0)] : $unsigned(reg179)))},
                  {({(~|reg172), (|forvar173)} ?
                          ((reg182 ^~ reg178) ~^ {wire165}) : {(reg174 && reg175)})}};
              reg183 <= $unsigned(wire163[(4'he):(3'h6)]);
            end
        end
      if (wire161[(5'h14):(3'h6)])
        begin
          reg184 <= $signed(((~^((reg183 | wire164) * (reg172 ?
              reg183 : wire166))) ^~ $signed((7'h41))));
          for (forvar185 = (1'h0); (forvar185 < (1'h1)); forvar185 = (forvar185 + (1'h1)))
            begin
              reg186 <= ((reg182 ?
                  reg176 : $signed({wire163,
                      (wire165 || reg179)})) >>> (^(~^reg177)));
              reg187 <= (($signed(($unsigned(wire167) ?
                          wire161 : $unsigned(reg182))) ?
                      {forvar185[(4'h8):(3'h4)]} : $signed({$signed(reg186)})) ?
                  reg171 : $signed((~|({forvar170} ?
                      (~&reg176) : $signed(wire161)))));
              reg188 <= $signed($unsigned($signed(reg184)));
            end
          for (forvar189 = (1'h0); (forvar189 < (3'h4)); forvar189 = (forvar189 + (1'h1)))
            begin
              reg190 = {$signed((^((~^wire162) ?
                      (8'ha4) : ((8'ha8) | forvar173)))),
                  $unsigned($signed({((8'hb9) <<< (8'hba))}))};
              reg191 <= (8'hb4);
            end
          reg192 = wire168;
        end
      else
        begin
          reg184 = (~&(~^((reg191 ~^ $unsigned((8'hb4))) ?
              (reg191[(3'h4):(2'h3)] ?
                  (forvar170 ?
                      reg176 : forvar185) : reg187[(1'h1):(1'h0)]) : ($signed(forvar170) ~^ $signed(reg178)))));
          reg185 = $unsigned($unsigned((~|(wire166[(2'h2):(1'h1)] >>> $unsigned(forvar185)))));
          for (forvar186 = (1'h0); (forvar186 < (2'h3)); forvar186 = (forvar186 + (1'h1)))
            begin
              reg187 <= ($signed(wire165) ?
                  (~|wire166[(3'h4):(1'h0)]) : (~&$unsigned((~^(&(7'h40))))));
              reg188 <= ($signed((~|(forvar180 ?
                  (wire164 ? reg185 : reg179) : (forvar189 ?
                      reg176 : (8'hac))))) == ((&wire167[(3'h6):(3'h5)]) ?
                  $unsigned({forvar185}) : (~^{(8'ha9)})));
              reg189 <= (~($unsigned(forvar189[(3'h4):(1'h0)]) ?
                  (~^(wire165[(5'h10):(1'h1)] ?
                      (reg192 ? reg174 : (8'hb8)) : {wire164,
                          reg183})) : $unsigned((~wire165[(4'h9):(4'h9)]))));
              reg190 <= wire164;
            end
        end
    end
  assign wire193 = $unsigned((reg171[(1'h0):(1'h0)] ?
                       (wire164 >> $unsigned({(8'haf)})) : ($unsigned((8'h9c)) > $signed({(8'hb6)}))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module136
#( parameter param153 = ((~|((((8'hba) ? (8'hb0) : (8'ha2)) ? ((8'ha4) ? (8'hab) : (8'hb3)) : ((8'hb7) ? (8'hb4) : (8'hbd))) ? {((7'h42) == (8'hb8)), (8'haa)} : {(~^(8'ha9))})) * {(+((+(8'hb8)) ? ((7'h44) >>> (8'ha7)) : (|(8'hbf))))})
, parameter param154 = (param153 >> (^~(8'ha8))) )
(y, clk, wire140, wire139, wire138, wire137);
  output wire [(32'h79):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h15):(1'h0)] wire140;
  input wire [(4'hc):(1'h0)] wire139;
  input wire signed [(4'h8):(1'h0)] wire138;
  input wire [(5'h11):(1'h0)] wire137;
  reg signed [(5'h10):(1'h0)] reg152 = (1'h0);
  reg [(3'h6):(1'h0)] reg151 = (1'h0);
  wire signed [(4'he):(1'h0)] wire150;
  wire [(3'h7):(1'h0)] wire149;
  wire signed [(4'ha):(1'h0)] wire148;
  reg [(3'h6):(1'h0)] reg147 = (1'h0);
  reg [(3'h4):(1'h0)] reg146 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire145;
  wire [(5'h10):(1'h0)] wire144;
  wire signed [(3'h5):(1'h0)] wire143;
  wire [(3'h6):(1'h0)] wire142;
  wire signed [(5'h15):(1'h0)] wire141;
  assign y = {reg152,
                 reg151,
                 wire150,
                 wire149,
                 wire148,
                 reg147,
                 reg146,
                 wire145,
                 wire144,
                 wire143,
                 wire142,
                 wire141,
                 (1'h0)};
  assign wire141 = wire139;
  assign wire142 = ($signed(wire137[(3'h4):(1'h1)]) ?
                       {wire141[(3'h6):(3'h4)]} : wire138[(3'h6):(1'h1)]);
  assign wire143 = ({($signed((wire138 ? wire138 : wire141)) ?
                           $unsigned($signed((8'ha8))) : wire141[(4'hb):(4'h8)])} | {$unsigned(((~&wire140) ?
                           ((8'hb2) ?
                               (8'hbf) : wire141) : wire142[(3'h5):(3'h4)])),
                       ($unsigned($unsigned(wire138)) ?
                           wire138 : $unsigned((wire141 ?
                               wire137 : wire137)))});
  assign wire144 = (^~(7'h41));
  assign wire145 = wire141[(3'h6):(3'h5)];
  always
    @(posedge clk) begin
      reg146 = $signed(wire142[(3'h4):(2'h2)]);
      reg147 = wire145[(1'h0):(1'h0)];
    end
  assign wire148 = $signed((8'hb2));
  assign wire149 = (&$unsigned(((~^(wire142 > wire138)) <= wire141)));
  assign wire150 = ($unsigned((wire141 ?
                       (|(~^reg146)) : wire141)) && (wire139[(4'hb):(3'h7)] ?
                       $signed((&$unsigned(wire144))) : wire141[(4'hc):(3'h6)]));
  always
    @(posedge clk) begin
      reg151 = (($signed($signed(wire150[(4'hc):(2'h2)])) ?
          $unsigned(((wire144 ? wire138 : wire145) >= {(8'hb4),
              reg147})) : (~&$unsigned((wire140 | wire143)))) | wire142);
      reg152 <= wire138;
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module427  (y, clk, wire432, wire431, wire430, wire429, wire428);
  output wire [(32'h28):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire432;
  input wire signed [(5'h15):(1'h0)] wire431;
  input wire signed [(4'ha):(1'h0)] wire430;
  input wire [(4'he):(1'h0)] wire429;
  input wire [(3'h7):(1'h0)] wire428;
  wire signed [(3'h7):(1'h0)] wire437;
  wire signed [(4'h8):(1'h0)] wire436;
  wire signed [(4'hb):(1'h0)] wire435;
  reg [(4'h9):(1'h0)] reg434 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg433 = (1'h0);
  assign y = {wire437, wire436, wire435, reg434, reg433, (1'h0)};
  always
    @(posedge clk) begin
      reg433 <= $signed(wire429);
      reg434 <= (~|$signed(wire431));
    end
  assign wire435 = wire431[(4'hb):(4'ha)];
  assign wire436 = wire428[(1'h0):(1'h0)];
  assign wire437 = wire429[(1'h0):(1'h0)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module254
#( parameter param418 = ((((((8'hb7) ? (8'hac) : (8'ha1)) && ((7'h44) > (8'hb4))) & {(~^(8'ha0)), (!(8'ha2))}) << (({(8'h9d), (8'h9e)} ? ((7'h40) >> (8'ha1)) : {(8'hb7), (8'hb0)}) ? (~|(+(8'hb9))) : (8'hb7))) ? (({((8'ha3) ? (8'hbf) : (8'hb6))} == ((8'hbb) ? (~&(8'hb8)) : (+(8'haf)))) | (((&(8'hbd)) ^ ((7'h40) ^ (8'h9e))) <= (8'h9f))) : {{(((8'ha3) >> (8'ha8)) ~^ ((8'hba) ? (8'ha1) : (7'h43)))}, ({((8'ha0) ? (8'ha1) : (8'h9f))} << ({(8'hb3)} ? ((8'ha5) ? (8'had) : (8'hb5)) : (8'hbf)))}) )
(y, clk, wire255, wire256, wire257, wire258);
  output wire [(32'h25c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire255;
  input wire signed [(4'hf):(1'h0)] wire256;
  input wire signed [(2'h3):(1'h0)] wire257;
  input wire signed [(5'h10):(1'h0)] wire258;
  wire signed [(3'h4):(1'h0)] wire417;
  wire [(4'hd):(1'h0)] wire416;
  reg [(4'ha):(1'h0)] reg415 = (1'h0);
  reg [(5'h10):(1'h0)] reg414 = (1'h0);
  reg [(4'hd):(1'h0)] reg413 = (1'h0);
  reg [(3'h7):(1'h0)] reg412 = (1'h0);
  reg [(5'h14):(1'h0)] reg411 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar410 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire409;
  wire [(4'hb):(1'h0)] wire408;
  wire [(4'hc):(1'h0)] wire259;
  reg [(5'h10):(1'h0)] reg260 = (1'h0);
  reg [(4'ha):(1'h0)] reg261 = (1'h0);
  reg [(5'h13):(1'h0)] reg262 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg263 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire264;
  wire [(3'h5):(1'h0)] wire265;
  wire [(4'he):(1'h0)] wire266;
  wire [(5'h11):(1'h0)] wire267;
  reg signed [(5'h11):(1'h0)] reg268 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar269 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg270 = (1'h0);
  reg [(3'h6):(1'h0)] forvar271 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg272 = (1'h0);
  reg [(3'h6):(1'h0)] reg273 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar274 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg275 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg276 = (1'h0);
  reg [(5'h12):(1'h0)] reg277 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg278 = (1'h0);
  reg [(5'h10):(1'h0)] reg279 = (1'h0);
  reg [(4'hf):(1'h0)] reg280 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar281 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg282 = (1'h0);
  reg [(3'h5):(1'h0)] reg283 = (1'h0);
  reg [(4'hd):(1'h0)] reg284 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg285 = (1'h0);
  reg [(4'ha):(1'h0)] reg286 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar287 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg288 = (1'h0);
  reg [(3'h6):(1'h0)] reg289 = (1'h0);
  reg [(2'h2):(1'h0)] reg290 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg291 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg292 = (1'h0);
  reg [(5'h13):(1'h0)] reg281 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire293;
  wire [(5'h10):(1'h0)] wire294;
  wire [(4'hd):(1'h0)] wire406;
  assign y = {wire417,
                 wire416,
                 reg415,
                 reg414,
                 reg413,
                 reg412,
                 reg411,
                 forvar410,
                 wire409,
                 wire408,
                 wire259,
                 reg260,
                 reg261,
                 reg262,
                 reg263,
                 wire264,
                 wire265,
                 wire266,
                 wire267,
                 reg268,
                 forvar269,
                 reg270,
                 forvar271,
                 reg272,
                 reg273,
                 forvar274,
                 reg275,
                 reg276,
                 reg277,
                 reg278,
                 reg279,
                 reg280,
                 forvar281,
                 reg282,
                 reg283,
                 reg284,
                 reg285,
                 reg286,
                 forvar287,
                 reg288,
                 reg289,
                 reg290,
                 reg291,
                 reg292,
                 reg281,
                 wire293,
                 wire294,
                 wire406,
                 (1'h0)};
  assign wire259 = $signed((!wire258));
  always
    @(posedge clk) begin
      reg260 <= (wire257 ?
          ($unsigned(wire256) ?
              (~&wire258) : wire258) : {wire258[(2'h2):(2'h2)]});
      reg261 <= (wire255 - $signed((($unsigned(reg260) < wire258) >> {(~wire258),
          (^reg260)})));
      reg262 = wire257[(2'h3):(2'h3)];
      reg263 <= $signed(((~reg262[(4'hb):(2'h2)]) <= {((reg261 ?
                  reg260 : wire257) ?
              $signed((8'haf)) : $unsigned((8'hb3)))}));
    end
  assign wire264 = ((~^reg261) ?
                       $unsigned(reg260[(2'h3):(1'h0)]) : $signed((8'hb6)));
  assign wire265 = wire257[(1'h1):(1'h0)];
  assign wire266 = reg260;
  assign wire267 = (wire255[(3'h4):(1'h1)] * wire264[(1'h1):(1'h1)]);
  always
    @(posedge clk) begin
      reg268 <= $signed(((^reg263[(4'hf):(4'h8)]) ?
          (wire257[(2'h3):(2'h3)] - $unsigned($unsigned(reg262))) : (reg261 <<< ({reg261} | reg260[(1'h1):(1'h0)]))));
      for (forvar269 = (1'h0); (forvar269 < (1'h1)); forvar269 = (forvar269 + (1'h1)))
        begin
          reg270 <= wire255;
          for (forvar271 = (1'h0); (forvar271 < (3'h4)); forvar271 = (forvar271 + (1'h1)))
            begin
              reg272 <= wire267;
            end
          reg273 <= ($signed((~|($unsigned(wire258) <<< (^~reg272)))) ?
              (8'hb8) : reg262[(4'hc):(4'ha)]);
        end
      for (forvar274 = (1'h0); (forvar274 < (2'h3)); forvar274 = (forvar274 + (1'h1)))
        begin
          reg275 <= (~((+(8'hbc)) ?
              $signed(wire267) : {(+$unsigned(wire265))}));
          reg276 <= (^~$unsigned(reg270));
          reg277 <= (~(((wire256[(4'ha):(4'h9)] != (reg260 ?
                  reg272 : (8'haf))) ?
              $signed({wire257}) : {reg273[(3'h5):(3'h5)],
                  $unsigned((8'hbf))}) || $unsigned($unsigned($signed(reg261)))));
          reg278 <= wire259;
          reg279 <= wire257;
        end
      reg280 <= ((|reg277[(4'hc):(3'h6)]) ?
          (~&(((~^wire255) ^~ (8'hbb)) | {{reg261},
              $signed(reg261)})) : wire258);
      if ((reg263 ? (8'hbd) : {(8'ha6)}))
        begin
          for (forvar281 = (1'h0); (forvar281 < (1'h1)); forvar281 = (forvar281 + (1'h1)))
            begin
              reg282 <= $signed($signed(((+(!reg260)) ?
                  ((reg263 <<< reg278) ?
                      (wire267 ?
                          forvar269 : wire255) : (~&reg261)) : ($signed(reg270) ?
                      $signed(reg280) : (wire257 ? reg262 : reg278)))));
              reg283 <= wire259[(2'h3):(2'h3)];
              reg284 <= $signed({({((8'h9f) <<< reg277)} | $unsigned($unsigned(reg283)))});
            end
          reg285 = $signed((7'h40));
          reg286 <= (forvar269[(4'hd):(4'h9)] + ({($unsigned(wire257) >>> forvar281),
                  reg285} ?
              $unsigned(reg280[(3'h7):(3'h6)]) : reg276[(4'ha):(3'h4)]));
          for (forvar287 = (1'h0); (forvar287 < (1'h0)); forvar287 = (forvar287 + (1'h1)))
            begin
              reg288 <= reg284;
              reg289 = $signed((~&$unsigned(({wire264} ?
                  reg268[(3'h4):(1'h1)] : reg275[(1'h1):(1'h1)]))));
              reg290 <= $unsigned(forvar269);
              reg291 = (8'hbc);
              reg292 <= (^wire265[(3'h4):(1'h1)]);
            end
        end
      else
        begin
          reg281 <= (!(^~((|{wire256, (8'hbe)}) ?
              ((reg285 > forvar287) ?
                  (reg275 >>> reg268) : {wire257}) : ((8'hb3) * $unsigned(reg283)))));
          reg282 <= ((~&$signed(((|(8'hb8)) ?
              $signed(forvar271) : $signed(reg277)))) >> $unsigned((|((~|wire266) ?
              $signed((8'hba)) : $unsigned(reg291)))));
          reg283 <= ((8'ha5) ?
              wire256[(4'hf):(4'h9)] : (forvar281 ?
                  {(reg291 >> wire257)} : {($signed(reg281) ?
                          $signed((8'hbb)) : (+reg279))}));
        end
    end
  assign wire293 = $signed((-$unsigned(reg273[(1'h1):(1'h1)])));
  assign wire294 = forvar269;
  module295 modinst407 (.wire296(reg261), .wire297(reg273), .wire299(wire264), .clk(clk), .wire300(wire258), .y(wire406), .wire298(reg272));
  assign wire408 = $signed(({(wire294 - reg276), wire264} ~^ {{(reg268 ?
                               (8'ha8) : reg291)}}));
  assign wire409 = {$unsigned(((+$signed(reg260)) ?
                           wire257[(1'h0):(1'h0)] : (wire406[(2'h3):(2'h2)] ?
                               (+wire258) : (forvar287 ? reg280 : wire266))))};
  always
    @(posedge clk) begin
      for (forvar410 = (1'h0); (forvar410 < (3'h4)); forvar410 = (forvar410 + (1'h1)))
        begin
          if ({(reg275[(2'h3):(2'h3)] ?
                  $unsigned($signed(reg272)) : (~|forvar281[(4'hc):(2'h3)])),
              reg286})
            begin
              reg411 <= $unsigned(reg270);
              reg412 <= reg276;
              reg413 <= (|{((~|(wire257 >>> reg286)) > ((wire256 ?
                      (8'ha1) : (8'hb3)) == reg276))});
              reg414 <= (wire259[(2'h3):(2'h2)] | wire255);
              reg415 <= reg273[(3'h5):(1'h1)];
            end
          else
            begin
              reg411 <= (((forvar410 <<< {(~|reg291),
                      (wire259 ?
                          wire264 : (8'hac))}) || reg415[(2'h3):(1'h1)]) ?
                  $unsigned(wire255[(1'h0):(1'h0)]) : ((~^$unsigned((reg280 * reg262))) ?
                      $unsigned(reg273) : (forvar410[(3'h6):(3'h6)] ?
                          $signed(reg278[(3'h7):(3'h5)]) : (reg280[(2'h3):(2'h2)] <= reg278))));
              reg412 = (($signed($signed((wire409 ? reg411 : forvar274))) ?
                      ((reg280[(2'h3):(1'h0)] ?
                          $unsigned((7'h40)) : {(8'h9c)}) ^ reg261[(4'ha):(2'h3)]) : {$unsigned(((8'hb1) ?
                              (7'h40) : reg277)),
                          reg411[(4'hf):(4'ha)]}) ?
                  forvar281 : (wire255 - (($signed(wire257) ?
                      $signed((8'hb0)) : wire265[(1'h0):(1'h0)]) > (^~$unsigned(reg412)))));
            end
        end
    end
  assign wire416 = $signed($signed(($signed((wire265 || reg282)) ?
                       $signed((wire293 > reg263)) : {(!reg412)})));
  assign wire417 = (reg263[(3'h6):(2'h3)] ?
                       $unsigned(wire408) : $signed(reg279[(2'h2):(1'h0)]));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module295
#( parameter param404 = ((!((8'hbb) ? ({(7'h44), (8'hbd)} << {(8'hbf)}) : {{(8'ha5), (8'hac)}})) <= {(7'h44), (~(|((8'haf) - (8'hb9))))})
, parameter param405 = ((((8'hb4) ? param404 : {(+param404)}) - ({(~&param404), {param404}} || ({param404} ? ((8'ha8) ? param404 : param404) : (^~(7'h41))))) > (&((param404 ? (8'hb6) : param404) ? (!{(8'ha4)}) : {(param404 ? param404 : param404)}))) )
(y, clk, wire300, wire299, wire298, wire297, wire296);
  output wire [(32'h2e4):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire300;
  input wire [(5'h10):(1'h0)] wire299;
  input wire signed [(4'h8):(1'h0)] wire298;
  input wire signed [(3'h6):(1'h0)] wire297;
  input wire [(4'ha):(1'h0)] wire296;
  reg [(5'h15):(1'h0)] reg403 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg402 = (1'h0);
  reg signed [(4'he):(1'h0)] reg401 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg400 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg399 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg398 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg397 = (1'h0);
  reg [(4'hf):(1'h0)] reg396 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg395 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg394 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar393 = (1'h0);
  reg [(4'hc):(1'h0)] reg392 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg391 = (1'h0);
  reg [(3'h6):(1'h0)] reg390 = (1'h0);
  reg [(2'h2):(1'h0)] reg389 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg388 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg387 = (1'h0);
  reg [(4'h9):(1'h0)] forvar382 = (1'h0);
  reg [(4'he):(1'h0)] reg381 = (1'h0);
  reg [(4'h9):(1'h0)] forvar380 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg386 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg385 = (1'h0);
  reg [(2'h2):(1'h0)] reg384 = (1'h0);
  reg [(3'h7):(1'h0)] reg383 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg382 = (1'h0);
  reg [(5'h12):(1'h0)] forvar381 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg380 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg379 = (1'h0);
  reg [(5'h12):(1'h0)] reg378 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg377 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg376 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar375 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire374;
  wire [(5'h12):(1'h0)] wire372;
  reg [(4'he):(1'h0)] reg324 = (1'h0);
  reg [(4'hd):(1'h0)] reg323 = (1'h0);
  reg [(2'h2):(1'h0)] reg322 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg321 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg320 = (1'h0);
  reg [(4'hd):(1'h0)] reg319 = (1'h0);
  reg [(5'h12):(1'h0)] reg318 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg317 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar316 = (1'h0);
  reg [(5'h14):(1'h0)] forvar315 = (1'h0);
  reg [(2'h3):(1'h0)] reg314 = (1'h0);
  reg [(4'hc):(1'h0)] reg313 = (1'h0);
  reg [(5'h11):(1'h0)] reg312 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg311 = (1'h0);
  reg [(3'h5):(1'h0)] reg310 = (1'h0);
  reg [(5'h12):(1'h0)] reg309 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar308 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar307 = (1'h0);
  reg [(5'h13):(1'h0)] reg306 = (1'h0);
  reg [(5'h14):(1'h0)] reg305 = (1'h0);
  reg [(4'he):(1'h0)] reg304 = (1'h0);
  reg [(5'h15):(1'h0)] reg303 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg302 = (1'h0);
  reg [(4'hf):(1'h0)] reg301 = (1'h0);
  assign y = {reg403,
                 reg402,
                 reg401,
                 reg400,
                 reg399,
                 reg398,
                 reg397,
                 reg396,
                 reg395,
                 reg394,
                 forvar393,
                 reg392,
                 reg391,
                 reg390,
                 reg389,
                 reg388,
                 reg387,
                 forvar382,
                 reg381,
                 forvar380,
                 reg386,
                 reg385,
                 reg384,
                 reg383,
                 reg382,
                 forvar381,
                 reg380,
                 reg379,
                 reg378,
                 reg377,
                 reg376,
                 forvar375,
                 wire374,
                 wire372,
                 reg324,
                 reg323,
                 reg322,
                 reg321,
                 reg320,
                 reg319,
                 reg318,
                 reg317,
                 forvar316,
                 forvar315,
                 reg314,
                 reg313,
                 reg312,
                 reg311,
                 reg310,
                 reg309,
                 forvar308,
                 forvar307,
                 reg306,
                 reg305,
                 reg304,
                 reg303,
                 reg302,
                 reg301,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg301 <= wire298[(1'h0):(1'h0)];
      reg302 <= reg301;
    end
  always
    @(posedge clk) begin
      reg303 <= $unsigned({$signed(((|wire298) ?
              (reg302 <<< wire298) : (wire299 >= wire299)))});
      reg304 <= {(wire298[(3'h6):(3'h5)] << ({$signed(wire299),
                  (wire296 ? reg303 : reg303)} ?
              ((wire296 ^~ reg302) ^~ (wire296 | (8'hb7))) : reg301)),
          ((({wire296, (8'hab)} ?
              (wire297 ?
                  (8'ha2) : reg303) : (^~(8'ha2))) * $unsigned($unsigned(wire297))) && reg302)};
      reg305 <= $signed(reg304[(4'he):(3'h6)]);
    end
  always
    @(posedge clk) begin
      reg306 <= reg305;
      for (forvar307 = (1'h0); (forvar307 < (2'h3)); forvar307 = (forvar307 + (1'h1)))
        begin
          for (forvar308 = (1'h0); (forvar308 < (2'h2)); forvar308 = (forvar308 + (1'h1)))
            begin
              reg309 <= $unsigned(($unsigned(((reg304 ^~ wire299) ^~ forvar308)) > ((reg305[(5'h13):(3'h6)] ?
                      $unsigned(reg305) : (reg303 ? wire299 : (8'hb4))) ?
                  (wire297 ?
                      (wire298 ? reg306 : reg304) : {wire298,
                          forvar307}) : $unsigned($unsigned(wire300)))));
              reg310 <= wire296;
              reg311 <= {reg302,
                  {reg301[(4'he):(4'hd)],
                      ({{reg304}} <= (~^((8'ha9) ~^ (8'ha6))))}};
              reg312 <= wire297;
            end
          reg313 <= $signed(reg304);
          reg314 <= reg301[(1'h1):(1'h1)];
        end
      for (forvar315 = (1'h0); (forvar315 < (3'h4)); forvar315 = (forvar315 + (1'h1)))
        begin
          for (forvar316 = (1'h0); (forvar316 < (2'h3)); forvar316 = (forvar316 + (1'h1)))
            begin
              reg317 = (^$unsigned($unsigned($signed(forvar315[(4'ha):(1'h1)]))));
              reg318 <= $unsigned($unsigned({((reg303 == reg309) < wire299[(3'h4):(3'h4)]),
                  (~&wire300[(4'h9):(1'h0)])}));
            end
          reg319 <= $unsigned($unsigned(reg314[(1'h1):(1'h0)]));
          reg320 = $signed(((forvar307 ?
                  wire298[(2'h3):(1'h0)] : (~|(reg305 ? forvar315 : (8'hac)))) ?
              reg311[(1'h0):(1'h0)] : {$signed(((8'hb3) ? (8'hb7) : reg313))}));
          reg321 <= $unsigned((reg304[(1'h1):(1'h0)] ?
              (((forvar308 ? reg304 : reg303) ?
                  (wire298 ^~ (8'hac)) : (reg317 >> wire299)) & $signed({(8'ha8)})) : ((|(|reg310)) ?
                  reg311 : reg319[(1'h1):(1'h1)])));
        end
    end
  always
    @(posedge clk) begin
      reg322 = wire298;
      reg323 = (^~((^wire297) ?
          $unsigned((8'ha4)) : ($signed($unsigned(wire296)) ~^ ($unsigned(wire299) >= (|reg318)))));
    end
  always
    @(posedge clk) begin
      reg324 <= forvar307[(1'h0):(1'h0)];
    end
  module325 modinst373 (.y(wire372), .wire327(reg313), .wire328(reg324), .wire326(reg304), .clk(clk), .wire329(forvar307));
  assign wire374 = $signed(((~&$unsigned(reg301)) <= reg319));
  always
    @(posedge clk) begin
      for (forvar375 = (1'h0); (forvar375 < (2'h2)); forvar375 = (forvar375 + (1'h1)))
        begin
          reg376 <= $signed(wire299);
          reg377 <= {$unsigned((~&$unsigned(forvar315[(4'ha):(3'h6)])))};
          reg378 <= ((~^(reg312[(4'hb):(3'h5)] == (reg376[(3'h7):(3'h7)] ?
                  $unsigned((7'h44)) : (!reg376)))) ?
              reg319 : forvar307[(2'h3):(1'h1)]);
          reg379 <= wire297[(3'h6):(1'h1)];
        end
      if (wire299)
        begin
          reg380 = wire374;
          for (forvar381 = (1'h0); (forvar381 < (2'h3)); forvar381 = (forvar381 + (1'h1)))
            begin
              reg382 = (~^reg321);
              reg383 <= $unsigned(reg382[(3'h4):(2'h3)]);
              reg384 <= reg380[(5'h11):(2'h3)];
              reg385 <= $unsigned(({(reg382[(2'h3):(1'h0)] - $unsigned(forvar316))} ~^ {(((8'ha3) ?
                      reg304 : reg322) > (^~reg324))}));
              reg386 <= {$unsigned($signed(reg323))};
            end
        end
      else
        begin
          for (forvar380 = (1'h0); (forvar380 < (1'h0)); forvar380 = (forvar380 + (1'h1)))
            begin
              reg381 <= reg317;
            end
          for (forvar382 = (1'h0); (forvar382 < (1'h1)); forvar382 = (forvar382 + (1'h1)))
            begin
              reg383 = wire372[(2'h2):(1'h0)];
              reg384 <= (~^wire299[(4'hc):(4'hb)]);
              reg385 <= ($unsigned(((+(reg385 ?
                      forvar308 : reg312)) >> $unsigned(forvar316))) ?
                  (&(wire372 || ((forvar308 ? reg380 : reg380) ?
                      (|reg318) : wire374[(4'h8):(3'h5)]))) : ($unsigned((!(wire298 ?
                          reg304 : reg379))) ?
                      ((~&forvar382[(3'h5):(2'h3)]) >>> (&$unsigned(forvar380))) : (|wire300[(2'h2):(1'h0)])));
              reg386 <= {{$signed((reg303 > (~wire300))),
                      (reg302 ?
                          (^~{wire374}) : ($unsigned(forvar308) && $signed(reg383)))}};
              reg387 <= $signed(($signed(((forvar316 ? wire297 : reg305) ?
                  $unsigned(reg381) : {forvar375})) && (+$unsigned((!reg324)))));
            end
          reg388 = $unsigned({($unsigned(wire297) < (~&$unsigned(reg320))),
              ({$signed(forvar315)} ?
                  ((reg302 ? reg387 : reg302) ?
                      reg323 : reg381[(4'hb):(4'hb)]) : (reg387 == (wire299 ^~ (8'hba))))});
          reg389 <= wire296;
          reg390 <= reg387[(4'h8):(4'h8)];
        end
      reg391 <= $signed(($unsigned((-reg386[(4'hc):(3'h5)])) < $signed((8'h9d))));
    end
  always
    @(posedge clk) begin
      reg392 <= $unsigned($unsigned(reg384[(2'h2):(2'h2)]));
      for (forvar393 = (1'h0); (forvar393 < (1'h1)); forvar393 = (forvar393 + (1'h1)))
        begin
          reg394 <= $signed($unsigned({({(8'hae),
                  reg392} ^ (forvar316 != reg390)),
              (^(8'ha2))}));
          reg395 = wire372[(5'h11):(2'h2)];
          reg396 <= $unsigned($unsigned(wire374[(4'h8):(1'h0)]));
          reg397 = (wire374 ?
              (reg396[(4'hc):(4'h9)] & ($signed({(8'hb6)}) && reg322)) : reg322);
        end
      reg398 <= ((!(+$unsigned(reg397))) | wire296);
    end
  always
    @(posedge clk) begin
      reg399 <= ($signed((reg323 || $signed($unsigned(reg320)))) ?
          $unsigned((^~$signed((~|(8'hbf))))) : forvar382);
      reg400 <= (-reg382);
      reg401 <= $signed($signed((&reg380)));
      reg402 <= $signed(reg378);
      reg403 <= forvar316[(1'h1):(1'h1)];
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module325  (y, clk, wire329, wire328, wire327, wire326);
  output wire [(32'h1de):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h3):(1'h0)] wire329;
  input wire [(4'he):(1'h0)] wire328;
  input wire [(4'hc):(1'h0)] wire327;
  input wire [(3'h6):(1'h0)] wire326;
  wire [(4'hd):(1'h0)] wire371;
  reg signed [(4'h8):(1'h0)] reg370 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg369 = (1'h0);
  reg [(5'h14):(1'h0)] reg368 = (1'h0);
  reg [(5'h15):(1'h0)] reg367 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire366;
  wire signed [(5'h10):(1'h0)] wire365;
  reg [(4'hb):(1'h0)] reg364 = (1'h0);
  reg [(4'he):(1'h0)] reg363 = (1'h0);
  wire [(4'hb):(1'h0)] wire362;
  wire signed [(5'h10):(1'h0)] wire361;
  wire signed [(4'ha):(1'h0)] wire360;
  wire signed [(5'h12):(1'h0)] wire359;
  reg [(2'h2):(1'h0)] reg358 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg357 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg356 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg355 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg354 = (1'h0);
  reg [(3'h5):(1'h0)] forvar353 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg352 = (1'h0);
  reg [(4'ha):(1'h0)] reg351 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg350 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg349 = (1'h0);
  reg [(5'h12):(1'h0)] reg348 = (1'h0);
  reg [(5'h15):(1'h0)] reg347 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg346 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg345 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg344 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg343 = (1'h0);
  reg [(3'h5):(1'h0)] reg342 = (1'h0);
  reg [(5'h11):(1'h0)] reg341 = (1'h0);
  reg [(2'h2):(1'h0)] reg340 = (1'h0);
  reg [(4'ha):(1'h0)] reg339 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar338 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg337 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg336 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg335 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg334 = (1'h0);
  reg [(2'h2):(1'h0)] forvar333 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg332 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg331 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg330 = (1'h0);
  assign y = {wire371,
                 reg370,
                 reg369,
                 reg368,
                 reg367,
                 wire366,
                 wire365,
                 reg364,
                 reg363,
                 wire362,
                 wire361,
                 wire360,
                 wire359,
                 reg358,
                 reg357,
                 reg356,
                 reg355,
                 reg354,
                 forvar353,
                 reg352,
                 reg351,
                 reg350,
                 reg349,
                 reg348,
                 reg347,
                 reg346,
                 reg345,
                 reg344,
                 reg343,
                 reg342,
                 reg341,
                 reg340,
                 reg339,
                 forvar338,
                 reg337,
                 reg336,
                 reg335,
                 reg334,
                 forvar333,
                 reg332,
                 reg331,
                 reg330,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg330 <= wire327[(3'h7):(3'h4)];
      reg331 <= ((($signed((!wire328)) ?
              {$signed((8'hb3))} : ((-reg330) * (wire328 * wire329))) >= wire329) ?
          $signed((+($unsigned(reg330) ?
              $unsigned(reg330) : (reg330 + wire328)))) : wire327);
      if ($signed($unsigned((^~(8'ha8)))))
        begin
          reg332 <= $signed($signed($unsigned(reg330)));
        end
      else
        begin
          reg332 <= (((((~&wire329) ^ (wire326 >>> wire329)) ~^ ((wire327 ?
                  wire326 : wire326) + {wire329,
                  reg331})) <= $signed((-$unsigned(wire326)))) ?
              $signed((^((reg332 * wire327) ?
                  {wire326, reg332} : {wire327,
                      (8'hb9)}))) : {wire327[(4'hc):(3'h4)]});
          for (forvar333 = (1'h0); (forvar333 < (1'h1)); forvar333 = (forvar333 + (1'h1)))
            begin
              reg334 = $signed((reg330[(2'h2):(1'h0)] ?
                  {forvar333, reg331[(4'ha):(3'h4)]} : ((wire328 ?
                      {wire328} : {wire326, (8'ha0)}) <= ((wire329 ?
                          (7'h44) : wire329) ?
                      $signed(reg331) : reg331[(2'h3):(2'h3)]))));
              reg335 <= (8'hac);
              reg336 <= ((|wire326) ? reg332 : reg331[(5'h12):(5'h11)]);
            end
          reg337 <= $signed($unsigned($unsigned({{wire326, wire327},
              (reg332 ? reg331 : wire327)})));
          for (forvar338 = (1'h0); (forvar338 < (2'h2)); forvar338 = (forvar338 + (1'h1)))
            begin
              reg339 <= {(wire326 ?
                      $signed({(reg334 ?
                              (8'hb4) : (8'hbd))}) : ((reg335[(1'h0):(1'h0)] ?
                          $unsigned(wire326) : (reg330 ?
                              reg334 : reg331)) || (forvar338 >>> $signed(reg332))))};
              reg340 <= $unsigned({((forvar333[(2'h2):(1'h1)] ?
                      (reg334 >> wire328) : (!(8'hb9))) - $unsigned($signed(wire329))),
                  ((8'ha2) && {(-wire329), (wire326 < reg336)})});
              reg341 <= reg335;
              reg342 <= ($signed(reg340) && (reg335[(2'h3):(2'h2)] ?
                  {$unsigned($unsigned(reg332))} : reg339));
            end
        end
      reg343 = (wire326[(1'h1):(1'h1)] ?
          (^$unsigned({forvar333,
              ((8'hbe) | reg331)})) : $signed(reg336[(4'h8):(1'h0)]));
    end
  always
    @(posedge clk) begin
      reg344 <= reg341;
      reg345 <= ({$unsigned(reg337)} ?
          $signed(((^{reg332, wire327}) ?
              $signed(reg330) : ((^~(8'haa)) ?
                  $signed(reg343) : (&reg332)))) : reg337[(3'h5):(3'h5)]);
      reg346 <= ($signed((reg339 - $signed((wire327 ? reg334 : wire327)))) ?
          forvar338 : reg336);
      reg347 = wire329;
      reg348 <= (reg336 * reg335[(3'h7):(3'h4)]);
    end
  always
    @(posedge clk) begin
      reg349 <= $signed(reg341[(1'h1):(1'h0)]);
      reg350 = {(8'hb4), $unsigned(($unsigned((~reg331)) >= (~&(-(8'hbb)))))};
    end
  always
    @(posedge clk) begin
      reg351 <= {$unsigned(({(|reg345),
              (wire326 ? reg342 : reg336)} << (8'hbd)))};
    end
  always
    @(posedge clk) begin
      reg352 <= $unsigned($signed((({reg334, (7'h40)} > (8'hb6)) < reg344)));
      for (forvar353 = (1'h0); (forvar353 < (1'h0)); forvar353 = (forvar353 + (1'h1)))
        begin
          reg354 <= reg334[(1'h1):(1'h1)];
          reg355 = (^((~(^~$unsigned(reg343))) ?
              (({wire326, reg351} ?
                  (reg342 ?
                      reg339 : reg340) : (~wire329)) || forvar333[(1'h1):(1'h0)]) : (wire327 > (8'ha6))));
          reg356 <= ((!$signed((|$signed(wire329)))) ?
              ((reg355 ?
                  forvar353[(3'h5):(1'h1)] : $signed(forvar353)) >>> ((8'h9f) >= (^~reg345))) : $signed(($signed($unsigned(reg349)) < $signed((8'h9d)))));
          reg357 = $signed(reg344);
          reg358 = $unsigned($unsigned((($signed(reg340) && ((8'hae) ?
                  reg356 : reg342)) ?
              wire329[(2'h3):(2'h2)] : (^reg335))));
        end
    end
  assign wire359 = (~&{reg342[(1'h1):(1'h1)]});
  assign wire360 = ((^((8'hb7) ?
                           reg331[(2'h3):(2'h3)] : reg355[(4'h8):(1'h1)])) ?
                       (^~($unsigned((^~reg334)) < (~{wire329}))) : {reg350,
                           ($unsigned((!(7'h42))) ?
                               ((-reg357) ?
                                   reg339 : {reg331,
                                       reg351}) : (reg344[(4'he):(3'h7)] << (^~reg351)))});
  assign wire361 = reg354[(1'h0):(1'h0)];
  assign wire362 = (reg332 ? (~|forvar353) : reg346[(1'h0):(1'h0)]);
  always
    @(posedge clk) begin
      reg363 <= ((((reg350 >= ((8'hae) ? wire327 : reg330)) ?
          reg332[(4'he):(2'h2)] : ((~|forvar333) ?
              (~^wire360) : (|wire362))) != (~^((reg351 < (8'ha4)) ?
          (reg340 <= forvar333) : $unsigned((8'h9c))))) && forvar338);
      reg364 <= (~|wire329[(2'h2):(1'h0)]);
    end
  assign wire365 = $signed(wire329);
  assign wire366 = ((^$unsigned(reg334)) ?
                       (&(~&(+wire326[(1'h0):(1'h0)]))) : $signed(($unsigned((8'hb5)) && {(wire362 ^ forvar353)})));
  always
    @(posedge clk) begin
      reg367 <= forvar353[(1'h0):(1'h0)];
      reg368 = ((&(reg344 ?
              $unsigned($signed(reg348)) : wire360[(1'h1):(1'h0)])) ?
          $unsigned(reg354) : ($signed((reg348[(1'h1):(1'h0)] <<< $signed(wire327))) << ($unsigned(reg356[(1'h0):(1'h0)]) > {$unsigned(reg351)})));
      reg369 <= (~^reg334);
      reg370 <= $signed(($signed((!$unsigned((8'ha7)))) ?
          reg337[(3'h5):(3'h5)] : (reg357[(2'h3):(1'h1)] << $signed(((8'ha9) ?
              wire365 : reg343)))));
    end
  assign wire371 = $unsigned($signed($unsigned(wire362)));
endmodule