(* use_dsp48="no" *) (* use_dsp="no" *) module top
#( parameter param290 = (~^({(~(~&(8'hb8)))} != ((!((8'hb0) * (8'hb9))) ? (((7'h44) ? (8'hbe) : (8'hb7)) >>> (8'ha8)) : ((+(8'hb6)) | ((8'hbe) ? (8'ha2) : (8'haf))))))
, parameter param291 = {((~|{(~(8'hba))}) ? (({param290} - (param290 ? param290 : param290)) || param290) : param290)} )
(y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h3ed):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire4;
  input wire [(2'h2):(1'h0)] wire3;
  input wire signed [(3'h5):(1'h0)] wire2;
  input wire signed [(4'ha):(1'h0)] wire1;
  input wire [(5'h14):(1'h0)] wire0;
  wire signed [(5'h12):(1'h0)] wire289;
  reg signed [(3'h5):(1'h0)] reg288 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg287 = (1'h0);
  reg [(4'hd):(1'h0)] reg286 = (1'h0);
  reg [(4'ha):(1'h0)] reg285 = (1'h0);
  reg [(2'h3):(1'h0)] reg284 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg283 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg282 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg281 = (1'h0);
  wire [(5'h13):(1'h0)] wire280;
  wire signed [(5'h12):(1'h0)] wire279;
  reg signed [(4'hc):(1'h0)] reg278 = (1'h0);
  reg [(4'hb):(1'h0)] reg277 = (1'h0);
  reg [(5'h14):(1'h0)] reg276 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg275 = (1'h0);
  reg [(2'h2):(1'h0)] reg274 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg273 = (1'h0);
  reg [(3'h4):(1'h0)] forvar272 = (1'h0);
  reg [(4'hf):(1'h0)] reg271 = (1'h0);
  reg [(3'h5):(1'h0)] reg270 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg269 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar268 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg267 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg266 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg265 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg264 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar263 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg262 = (1'h0);
  reg [(5'h10):(1'h0)] reg261 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg260 = (1'h0);
  wire [(5'h11):(1'h0)] wire259;
  wire signed [(5'h11):(1'h0)] wire258;
  reg [(4'hd):(1'h0)] reg257 = (1'h0);
  reg signed [(4'he):(1'h0)] reg256 = (1'h0);
  reg [(4'hc):(1'h0)] reg255 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg254 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg253 = (1'h0);
  reg [(5'h13):(1'h0)] reg252 = (1'h0);
  reg [(3'h4):(1'h0)] reg251 = (1'h0);
  reg [(4'ha):(1'h0)] reg250 = (1'h0);
  reg [(4'h8):(1'h0)] reg249 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg248 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar247 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg246 = (1'h0);
  reg [(4'h9):(1'h0)] reg245 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg244 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg243 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar242 = (1'h0);
  reg [(4'hc):(1'h0)] reg241 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg240 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar239 = (1'h0);
  reg [(2'h2):(1'h0)] reg238 = (1'h0);
  reg [(3'h7):(1'h0)] reg237 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg236 = (1'h0);
  reg [(4'hf):(1'h0)] reg235 = (1'h0);
  reg [(3'h6):(1'h0)] reg234 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire233;
  wire signed [(4'hd):(1'h0)] wire207;
  wire signed [(4'hf):(1'h0)] wire159;
  wire [(3'h7):(1'h0)] wire157;
  wire [(5'h13):(1'h0)] wire30;
  reg signed [(4'hd):(1'h0)] reg29 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg28 = (1'h0);
  reg [(4'hb):(1'h0)] reg27 = (1'h0);
  reg [(5'h15):(1'h0)] reg26 = (1'h0);
  reg [(5'h10):(1'h0)] reg25 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg24 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg23 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg22 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar21 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar20 = (1'h0);
  reg [(5'h10):(1'h0)] reg19 = (1'h0);
  reg [(4'h8):(1'h0)] reg18 = (1'h0);
  reg [(4'hc):(1'h0)] reg17 = (1'h0);
  reg [(2'h2):(1'h0)] reg16 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg15 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg14 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg13 = (1'h0);
  reg signed [(4'he):(1'h0)] reg12 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg11 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg10 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg9 = (1'h0);
  reg [(2'h3):(1'h0)] forvar8 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar7 = (1'h0);
  reg [(4'hf):(1'h0)] reg6 = (1'h0);
  wire [(3'h6):(1'h0)] wire5;
  wire [(2'h3):(1'h0)] wire231;
  assign y = {wire289,
                 reg288,
                 reg287,
                 reg286,
                 reg285,
                 reg284,
                 reg283,
                 reg282,
                 reg281,
                 wire280,
                 wire279,
                 reg278,
                 reg277,
                 reg276,
                 reg275,
                 reg274,
                 reg273,
                 forvar272,
                 reg271,
                 reg270,
                 reg269,
                 forvar268,
                 reg267,
                 reg266,
                 reg265,
                 reg264,
                 forvar263,
                 reg262,
                 reg261,
                 reg260,
                 wire259,
                 wire258,
                 reg257,
                 reg256,
                 reg255,
                 reg254,
                 reg253,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 reg248,
                 forvar247,
                 reg246,
                 reg245,
                 reg244,
                 reg243,
                 forvar242,
                 reg241,
                 reg240,
                 forvar239,
                 reg238,
                 reg237,
                 reg236,
                 reg235,
                 reg234,
                 wire233,
                 wire207,
                 wire159,
                 wire157,
                 wire30,
                 reg29,
                 reg28,
                 reg27,
                 reg26,
                 reg25,
                 reg24,
                 reg23,
                 reg22,
                 forvar21,
                 forvar20,
                 reg19,
                 reg18,
                 reg17,
                 reg16,
                 reg15,
                 reg14,
                 reg13,
                 reg12,
                 reg11,
                 reg10,
                 reg9,
                 forvar8,
                 forvar7,
                 reg6,
                 wire5,
                 wire231,
                 (1'h0)};
  assign wire5 = wire4[(3'h4):(1'h0)];
  always
    @(posedge clk) begin
      reg6 <= $signed(wire0[(5'h13):(2'h3)]);
      for (forvar7 = (1'h0); (forvar7 < (1'h1)); forvar7 = (forvar7 + (1'h1)))
        begin
          for (forvar8 = (1'h0); (forvar8 < (2'h3)); forvar8 = (forvar8 + (1'h1)))
            begin
              reg9 <= $signed(wire4);
              reg10 <= {wire0};
              reg11 <= {$signed(wire4)};
              reg12 <= (wire0[(3'h6):(2'h2)] ?
                  ($signed($signed(wire2)) * wire3) : (!(8'hb9)));
              reg13 = ({(((reg10 || forvar7) + $unsigned(reg11)) ?
                      ((wire5 ^ wire3) != $signed(reg12)) : ({wire2, (8'hbd)} ?
                          reg6 : wire4[(3'h6):(3'h4)]))} ^~ (^~({$signed(wire3)} > (8'haa))));
            end
          reg14 <= reg6[(4'h8):(2'h3)];
          reg15 = (+$signed($unsigned(reg13)));
          reg16 <= {$unsigned({(-reg6[(3'h5):(2'h3)])})};
        end
      reg17 <= (~^wire0[(4'hc):(1'h1)]);
      reg18 <= wire3[(1'h0):(1'h0)];
      reg19 <= $signed((((~reg15[(1'h1):(1'h0)]) < ({reg18,
              reg9} << $signed(reg16))) ?
          (~&(reg6[(4'hd):(4'h8)] && (^reg12))) : $unsigned({(^~reg15),
              {(8'hbe)}})));
    end
  always
    @(posedge clk) begin
      for (forvar20 = (1'h0); (forvar20 < (2'h2)); forvar20 = (forvar20 + (1'h1)))
        begin
          for (forvar21 = (1'h0); (forvar21 < (2'h3)); forvar21 = (forvar21 + (1'h1)))
            begin
              reg22 <= reg10;
              reg23 <= (~^$unsigned((((reg6 ? wire0 : reg13) != (~^reg9)) ?
                  (&((8'hbe) >>> reg22)) : wire1[(4'h9):(3'h5)])));
              reg24 = (&wire1);
            end
          reg25 <= $signed({($unsigned($signed(forvar7)) ^~ reg17),
              (forvar20 ?
                  (wire4[(3'h5):(3'h5)] ?
                      (reg17 + reg16) : (wire1 >> reg19)) : (^forvar7))});
          reg26 = {(~^(!(~|{reg11})))};
        end
      reg27 <= (-(&(wire2 && reg18)));
      reg28 = (reg14 ? (-forvar8) : ($signed($signed((~^(7'h43)))) ^ wire2));
      reg29 <= (!$signed($unsigned((8'hb0))));
    end
  assign wire30 = wire5;
  module31 modinst158 (.clk(clk), .y(wire157), .wire33(reg17), .wire35(reg10), .wire34(reg27), .wire32(reg11));
  assign wire159 = (8'ha9);
  module160 modinst208 (.wire165(wire4), .clk(clk), .wire163(reg17), .wire164(reg25), .wire161(reg19), .wire162(reg14), .y(wire207));
  module209 modinst232 (.wire210(reg27), .wire214(reg13), .wire213(reg17), .y(wire231), .wire211(reg15), .clk(clk), .wire212(reg14));
  assign wire233 = {{{(!{reg16})}, $unsigned(reg29[(4'ha):(3'h5)])}};
  always
    @(posedge clk) begin
      reg234 <= reg23;
    end
  always
    @(posedge clk) begin
      reg235 <= (8'hbd);
      reg236 = (((reg12[(1'h0):(1'h0)] ?
          (~&$unsigned(reg26)) : ($signed((8'hb8)) ^ (8'had))) ^~ (reg17[(4'hb):(3'h7)] ?
          $unsigned({reg22, reg25}) : ({reg15} ?
              $signed(reg26) : (wire1 << (8'hbc))))) && forvar20[(2'h2):(2'h2)]);
      reg237 <= wire4[(5'h12):(3'h7)];
      reg238 = (wire207 ?
          ((+wire157[(2'h3):(1'h1)]) || (reg235[(1'h1):(1'h1)] | (+$unsigned((8'hbe))))) : (((~^((8'ha8) ?
                      reg235 : reg235)) ?
                  $unsigned($signed(forvar21)) : (-reg15)) ?
              ((^~(-(8'haa))) < ((~forvar8) | reg14[(4'hf):(4'hc)])) : ($signed((reg29 != reg14)) >> wire5)));
      for (forvar239 = (1'h0); (forvar239 < (2'h2)); forvar239 = (forvar239 + (1'h1)))
        begin
          reg240 <= wire2[(1'h1):(1'h1)];
          reg241 <= ({((wire30 ? reg23 : (wire233 << reg24)) || {(reg16 ?
                      reg12 : reg22),
                  wire233[(2'h2):(1'h0)]})} | (reg26 ?
              $unsigned((8'ha6)) : (($signed((8'had)) ?
                      $unsigned((8'ha4)) : reg28) ?
                  $unsigned(wire3[(2'h2):(2'h2)]) : (8'hb5))));
          for (forvar242 = (1'h0); (forvar242 < (2'h3)); forvar242 = (forvar242 + (1'h1)))
            begin
              reg243 <= {reg235[(3'h6):(2'h2)],
                  (wire4[(5'h12):(4'h8)] ?
                      $unsigned(({reg25} != $unsigned(reg236))) : forvar21)};
              reg244 <= (8'hab);
              reg245 = $unsigned({((~&wire1[(2'h3):(2'h3)]) ?
                      {reg16, forvar20} : $unsigned($signed(forvar239))),
                  reg11[(4'hd):(4'hb)]});
            end
          reg246 <= (wire1 > (^~$signed((~^$signed(reg17)))));
          for (forvar247 = (1'h0); (forvar247 < (1'h1)); forvar247 = (forvar247 + (1'h1)))
            begin
              reg248 = reg244[(1'h1):(1'h0)];
              reg249 <= {(~^((&(reg240 ? reg12 : reg17)) <= $signed(reg240)))};
              reg250 <= {$signed(({reg235} << $unsigned((reg6 ?
                      wire233 : wire1)))),
                  (+wire207[(1'h0):(1'h0)])};
              reg251 <= $signed((8'h9d));
              reg252 <= $signed((8'hb6));
            end
        end
    end
  always
    @(posedge clk) begin
      reg253 = forvar242[(1'h1):(1'h0)];
      reg254 = (({{(&(8'haa))},
          reg246[(4'ha):(4'ha)]} == ((forvar20[(3'h7):(3'h4)] ?
              forvar247 : forvar7[(1'h0):(1'h0)]) ?
          (!$signed((8'hbe))) : (~reg13[(2'h3):(2'h3)]))) >> $unsigned((wire159 && (~|{reg249,
          wire233}))));
      reg255 <= ($signed(forvar242) ?
          $unsigned({($unsigned(reg26) ?
                  (~(8'hb4)) : (forvar21 != reg14))}) : $signed($unsigned(reg9)));
      reg256 = (~|(^~$unsigned((reg240[(2'h3):(1'h0)] >>> $signed(reg29)))));
      reg257 <= reg28[(2'h2):(1'h0)];
    end
  assign wire258 = reg238[(1'h1):(1'h1)];
  assign wire259 = ({(!(8'hb7))} * ($signed($signed((8'h9d))) ?
                       (~^wire231) : ({(reg253 ~^ reg24)} <= forvar7)));
  always
    @(posedge clk) begin
      reg260 <= $signed(({$unsigned($unsigned(wire3)),
              (^~wire0[(4'hd):(4'hd)])} ?
          reg25[(3'h6):(2'h2)] : reg27));
      reg261 <= $signed($signed($unsigned((~^$signed(reg256)))));
    end
  always
    @(posedge clk) begin
      reg262 <= $unsigned({reg9[(4'hd):(3'h6)]});
      for (forvar263 = (1'h0); (forvar263 < (1'h0)); forvar263 = (forvar263 + (1'h1)))
        begin
          reg264 <= $unsigned(reg248[(2'h2):(2'h2)]);
          reg265 <= ($unsigned($signed((-((8'hb6) ?
              reg22 : reg28)))) >>> ((~^((reg240 ? reg248 : reg245) ?
                  (~&(8'hb1)) : $unsigned((8'hb7)))) ?
              $unsigned($unsigned(forvar8[(2'h2):(1'h1)])) : (^(!(wire3 < wire233)))));
          reg266 <= (reg235[(4'h8):(3'h6)] ?
              $unsigned($signed(((^~wire4) != $signed(reg19)))) : reg248[(1'h0):(1'h0)]);
          reg267 <= ((~{({reg251, reg25} + reg251),
              (reg9[(4'ha):(1'h1)] & reg10[(3'h6):(2'h2)])}) <= reg25);
          for (forvar268 = (1'h0); (forvar268 < (1'h1)); forvar268 = (forvar268 + (1'h1)))
            begin
              reg269 = (({$signed((-(8'ha3))),
                      $unsigned((~forvar21))} | ({(wire159 ?
                              reg23 : forvar20)} ?
                      ((~reg255) ^ $unsigned(reg17)) : $signed($signed((8'haf))))) ?
                  (!$unsigned(forvar247)) : wire5[(3'h4):(2'h2)]);
              reg270 <= wire157;
              reg271 <= reg249;
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar272 = (1'h0); (forvar272 < (1'h1)); forvar272 = (forvar272 + (1'h1)))
        begin
          reg273 <= (($signed(($unsigned(reg245) ^ $signed(wire231))) ?
              $unsigned({(reg27 <= (8'hb8)),
                  $unsigned(reg269)}) : reg12[(3'h4):(2'h2)]) || reg235[(4'hd):(2'h3)]);
          reg274 = $signed((8'h9d));
        end
      reg275 = (+$unsigned(reg249[(1'h1):(1'h0)]));
      reg276 <= {{(((reg19 ? (8'hba) : (8'hb5)) ?
                  {reg26, reg256} : ((8'h9c) ?
                      forvar20 : (8'hbf))) && ((reg273 ?
                  (8'hbd) : reg264) != reg270[(1'h1):(1'h1)])),
              $signed($unsigned($signed(forvar272)))}};
      reg277 <= (!reg238);
      reg278 <= reg17[(4'h8):(2'h3)];
    end
  assign wire279 = ((($unsigned($signed(forvar272)) ?
                           ((reg274 && (8'ha1)) + {(8'h9e),
                               forvar268}) : reg267[(3'h4):(2'h2)]) ?
                       {(wire159 << $unsigned(wire4))} : $signed($signed((reg271 ^~ reg278)))) << forvar247[(4'ha):(3'h6)]);
  assign wire280 = ($signed(reg6[(3'h4):(1'h1)]) > {(wire0 | (~^(~&reg246))),
                       ($unsigned((8'hbb)) ?
                           reg237 : $unsigned((wire233 ? reg241 : reg235)))});
  always
    @(posedge clk) begin
      reg281 <= (({((reg277 * (8'hbf)) ? (8'ha1) : {reg274, wire1}), reg18} ?
          (($signed(reg257) ?
              wire2[(2'h3):(2'h3)] : (8'h9e)) & $unsigned((reg277 ?
              reg260 : reg265))) : {(((8'ha0) ? reg16 : forvar239) ?
                  $unsigned(wire207) : reg278[(4'h8):(4'h8)]),
              ($unsigned(reg23) >> reg10[(2'h2):(1'h1)])}) ^ $signed(((&(-(8'hbf))) ?
          ((~reg266) ? (8'hac) : reg27) : reg10[(3'h6):(2'h2)])));
      reg282 = reg19[(3'h7):(3'h4)];
      reg283 <= {$signed(reg264[(1'h1):(1'h1)]),
          $unsigned($signed($signed(reg11[(1'h1):(1'h0)])))};
      reg284 <= reg17[(3'h6):(2'h2)];
      reg285 <= ($unsigned(wire4) ?
          ((7'h43) << (~^wire0)) : $unsigned(((reg255[(3'h6):(2'h3)] - wire279) ?
              (forvar263[(4'hf):(3'h6)] < reg266) : (wire159[(4'hb):(3'h4)] ?
                  $unsigned(reg270) : (reg12 ? reg284 : reg29)))));
    end
  always
    @(posedge clk) begin
      reg286 = (!(+((8'hb0) ?
          $unsigned((~reg248)) : ((reg278 ? reg22 : (8'hb2)) - (+reg13)))));
      reg287 = $signed((^~($signed($signed((8'had))) ?
          (~reg23[(4'hc):(3'h5)]) : $signed((+reg266)))));
      reg288 <= $unsigned(($unsigned((reg274 ?
              ((8'ha4) ? reg28 : wire157) : (reg255 >>> (8'hab)))) ?
          (~reg9) : wire157[(2'h2):(1'h0)]));
    end
  assign wire289 = $signed({(($unsigned((7'h40)) ?
                           $unsigned(reg285) : forvar263) ~^ reg285[(3'h4):(1'h0)])});
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module209
#( parameter param230 = {(((-((8'hb5) ^~ (8'hb0))) ? (7'h44) : (((8'hbf) ? (8'hb1) : (8'hab)) ^ ((8'hb1) ? (7'h40) : (7'h43)))) ? {{(^~(8'h9d)), ((8'hab) ? (8'hbd) : (8'h9d))}} : (~^(^~(-(8'hbd)))))} )
(y, clk, wire214, wire213, wire212, wire211, wire210);
  output wire [(32'hc6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire214;
  input wire [(4'ha):(1'h0)] wire213;
  input wire signed [(5'h11):(1'h0)] wire212;
  input wire signed [(3'h5):(1'h0)] wire211;
  input wire signed [(4'hb):(1'h0)] wire210;
  wire signed [(5'h10):(1'h0)] wire229;
  wire [(3'h7):(1'h0)] wire228;
  reg signed [(4'hb):(1'h0)] reg227 = (1'h0);
  wire [(5'h12):(1'h0)] wire226;
  wire [(3'h5):(1'h0)] wire225;
  wire [(2'h3):(1'h0)] wire224;
  reg [(5'h14):(1'h0)] reg223 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg222 = (1'h0);
  reg [(4'hc):(1'h0)] reg221 = (1'h0);
  reg [(4'h8):(1'h0)] reg220 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg219 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar218 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg217 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg216 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg215 = (1'h0);
  assign y = {wire229,
                 wire228,
                 reg227,
                 wire226,
                 wire225,
                 wire224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 reg219,
                 forvar218,
                 reg217,
                 reg216,
                 reg215,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg215 <= ($signed($unsigned({(&wire213)})) ?
          $signed(wire210) : (~^$signed(({wire211} ?
              $signed(wire210) : (^wire210)))));
      reg216 = (~|{(wire211[(2'h2):(1'h0)] & {(wire211 ~^ wire213)})});
      reg217 <= $signed(($signed(($signed(reg216) ?
              $signed(wire214) : (!wire212))) ?
          $signed(reg215) : $unsigned((~wire210[(4'h9):(3'h6)]))));
      for (forvar218 = (1'h0); (forvar218 < (2'h2)); forvar218 = (forvar218 + (1'h1)))
        begin
          reg219 <= reg216;
          reg220 <= ($unsigned(($unsigned({(8'hae),
                  (8'hb1)}) ^ (forvar218[(3'h6):(3'h6)] ?
                  wire212[(5'h10):(4'he)] : (~|wire212)))) ?
              {$signed($signed(wire213[(3'h6):(1'h1)]))} : $signed({reg217[(4'ha):(2'h2)],
                  ($signed(wire213) ? $signed(reg215) : $signed(reg219))}));
          reg221 <= ($unsigned($signed($signed($signed(wire211)))) ^ (+$signed((8'ha1))));
          reg222 <= $unsigned((8'h9c));
        end
      reg223 = $unsigned((($signed((|(8'hb2))) >= $unsigned((reg215 ?
          wire213 : reg221))) >>> $unsigned($signed((&(8'ha5))))));
    end
  assign wire224 = (wire212 >>> reg217[(3'h6):(1'h1)]);
  assign wire225 = (&{wire210[(1'h0):(1'h0)]});
  assign wire226 = (((reg220 ?
                           (+wire214) : {{wire210,
                                   reg221}}) == $unsigned(($signed(reg223) ^~ wire211[(2'h2):(2'h2)]))) ?
                       $unsigned($unsigned((forvar218[(4'ha):(1'h0)] | (-forvar218)))) : {reg221});
  always
    @(posedge clk) begin
      reg227 <= reg221[(4'hc):(4'ha)];
    end
  assign wire228 = (8'haa);
  assign wire229 = (^~reg223[(4'hf):(1'h0)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module160
#( parameter param206 = (({(+{(8'ha3), (8'hb3)})} ? ((((8'h9d) || (8'ha5)) ? (|(8'haf)) : ((8'haf) ? (8'hb2) : (8'hbc))) ? (+((8'hab) >= (8'hba))) : (~|((8'hb2) + (8'hb2)))) : (8'hab)) ? ((+{(|(7'h44)), (8'h9e)}) ? ((~&((8'had) ? (8'hab) : (8'ha6))) - {((8'ha2) || (8'ha6))}) : (^~(((8'ha9) <= (8'hb5)) != ((8'hac) <<< (8'ha4))))) : (((!(~|(7'h40))) + {((8'hb5) ? (8'haf) : (7'h44)), (^~(8'ha5))}) ? (~^{((8'ha2) <<< (7'h42)), ((8'hb0) ? (8'h9e) : (8'ha6))}) : (((^~(8'hb8)) ? {(8'ha4), (8'hac)} : ((8'hb0) * (8'hb9))) || (|{(8'ha9)})))) )
(y, clk, wire165, wire164, wire163, wire162, wire161);
  output wire [(32'h1b4):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire165;
  input wire [(4'hb):(1'h0)] wire164;
  input wire signed [(2'h2):(1'h0)] wire163;
  input wire signed [(4'he):(1'h0)] wire162;
  input wire [(5'h10):(1'h0)] wire161;
  reg signed [(4'h8):(1'h0)] reg205 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg204 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire203;
  wire signed [(2'h3):(1'h0)] wire202;
  reg signed [(5'h12):(1'h0)] reg201 = (1'h0);
  reg [(3'h6):(1'h0)] reg200 = (1'h0);
  reg [(4'ha):(1'h0)] reg199 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg198 = (1'h0);
  reg [(4'hf):(1'h0)] reg197 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar196 = (1'h0);
  reg [(4'h8):(1'h0)] reg195 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg194 = (1'h0);
  reg [(5'h13):(1'h0)] reg193 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg192 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg191 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg190 = (1'h0);
  reg [(4'hb):(1'h0)] forvar189 = (1'h0);
  reg [(3'h7):(1'h0)] forvar188 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg187 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg186 = (1'h0);
  reg [(4'h8):(1'h0)] reg185 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg184 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg183 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg182 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar181 = (1'h0);
  reg [(2'h2):(1'h0)] reg180 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg179 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg178 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar177 = (1'h0);
  reg [(3'h6):(1'h0)] reg176 = (1'h0);
  reg [(5'h13):(1'h0)] reg175 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar174 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg173 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire172;
  reg signed [(3'h6):(1'h0)] reg171 = (1'h0);
  reg signed [(4'he):(1'h0)] reg170 = (1'h0);
  reg [(4'ha):(1'h0)] reg169 = (1'h0);
  reg [(3'h7):(1'h0)] reg168 = (1'h0);
  reg [(4'hc):(1'h0)] reg167 = (1'h0);
  reg [(4'he):(1'h0)] reg166 = (1'h0);
  assign y = {reg205,
                 reg204,
                 wire203,
                 wire202,
                 reg201,
                 reg200,
                 reg199,
                 reg198,
                 reg197,
                 forvar196,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 reg191,
                 reg190,
                 forvar189,
                 forvar188,
                 reg187,
                 reg186,
                 reg185,
                 reg184,
                 reg183,
                 reg182,
                 forvar181,
                 reg180,
                 reg179,
                 reg178,
                 forvar177,
                 reg176,
                 reg175,
                 forvar174,
                 reg173,
                 wire172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg166 <= wire165[(1'h0):(1'h0)];
      reg167 <= wire163;
    end
  always
    @(posedge clk) begin
      reg168 <= {{(((wire163 >= wire163) + (wire165 != wire162)) == $signed(wire165)),
              wire161[(1'h0):(1'h0)]},
          ((8'hb2) <= ($signed($unsigned(reg167)) - ((8'h9f) ?
              (~|reg166) : (wire163 ? wire162 : wire163))))};
      reg169 = $unsigned($signed((-(+{wire164, (8'haa)}))));
      reg170 <= ((~wire162[(4'he):(4'hd)]) ?
          $signed(wire164) : {wire163[(1'h0):(1'h0)],
              $unsigned(reg167[(2'h3):(1'h1)])});
      reg171 <= ((!((((8'h9f) - reg166) ?
          {reg166} : reg166) && reg166[(4'he):(4'ha)])) <<< reg170[(2'h2):(1'h1)]);
    end
  assign wire172 = $signed(((~^($signed(reg168) ?
                           reg171[(3'h5):(1'h0)] : (reg167 ?
                               wire163 : wire164))) ?
                       (($unsigned((8'hbf)) & (reg171 ?
                           reg171 : wire161)) >= $signed((8'haf))) : $unsigned(wire164[(3'h4):(2'h2)])));
  always
    @(posedge clk) begin
      reg173 <= (((&(reg168[(3'h4):(2'h2)] ? wire172[(3'h6):(2'h3)] : reg166)) ?
          (^~(^{wire165,
              wire163})) : reg169) < (^$signed(wire164[(1'h1):(1'h0)])));
      for (forvar174 = (1'h0); (forvar174 < (2'h3)); forvar174 = (forvar174 + (1'h1)))
        begin
          reg175 <= ($signed((!{reg168})) ?
              wire164 : $unsigned((wire165[(1'h0):(1'h0)] ^~ (reg169[(2'h3):(2'h3)] - ((8'hbd) ?
                  wire172 : reg173)))));
          reg176 <= $signed({$signed(({(8'ha3), forvar174} ?
                  $signed(reg168) : reg173)),
              ($unsigned((reg171 ? reg168 : (8'haf))) * {reg168[(3'h7):(1'h1)],
                  (wire164 ^~ reg170)})});
          for (forvar177 = (1'h0); (forvar177 < (2'h2)); forvar177 = (forvar177 + (1'h1)))
            begin
              reg178 <= (($unsigned($signed({(8'hb3)})) <= (|$signed($signed(reg166)))) << $signed($unsigned({$unsigned(reg171),
                  {wire163, (8'ha6)}})));
            end
          reg179 = $signed(reg168);
          reg180 <= (($signed(($unsigned(reg171) ?
                  (|reg167) : {reg171, (8'ha6)})) ?
              $signed(reg170[(3'h6):(2'h3)]) : {wire165}) == reg167);
        end
      for (forvar181 = (1'h0); (forvar181 < (2'h2)); forvar181 = (forvar181 + (1'h1)))
        begin
          reg182 <= reg173[(4'h9):(1'h1)];
          reg183 <= forvar174[(2'h2):(2'h2)];
          reg184 <= (reg176 ?
              ({reg180, $signed($unsigned(reg179))} ?
                  $unsigned($unsigned(reg169[(3'h5):(1'h1)])) : reg173[(4'h8):(4'h8)]) : $unsigned(wire163));
          reg185 <= (&wire163[(1'h1):(1'h0)]);
          reg186 <= $unsigned((-(^(reg180 ?
              (reg176 ? (8'ha6) : forvar174) : $signed((7'h41))))));
        end
      reg187 = ((reg166[(4'ha):(3'h7)] ?
              wire161[(5'h10):(3'h5)] : (!reg186[(4'h9):(3'h6)])) ?
          reg175[(4'h8):(3'h6)] : {((~|(~&reg178)) ?
                  forvar174[(3'h6):(2'h3)] : reg168[(3'h5):(1'h1)])});
    end
  always
    @(posedge clk) begin
      for (forvar188 = (1'h0); (forvar188 < (3'h4)); forvar188 = (forvar188 + (1'h1)))
        begin
          for (forvar189 = (1'h0); (forvar189 < (3'h4)); forvar189 = (forvar189 + (1'h1)))
            begin
              reg190 <= $signed((forvar174 ?
                  (+$unsigned((^~reg176))) : (reg185[(3'h5):(3'h5)] ?
                      $signed(((7'h41) ? (8'hae) : forvar174)) : (reg184 ?
                          (~^wire161) : (~&reg178)))));
              reg191 = (forvar189[(1'h0):(1'h0)] ?
                  reg176 : ($unsigned(($signed(forvar189) ?
                          (~(8'h9e)) : $unsigned(reg170))) ?
                      ($signed((reg171 ?
                          (8'hae) : wire165)) - (((8'hbc) || reg173) ?
                          (wire161 ^~ reg170) : reg180)) : ((&(reg185 ?
                              (8'ha7) : reg169)) ?
                          reg167[(4'hb):(3'h4)] : reg180[(1'h0):(1'h0)])));
              reg192 <= (~&$signed($unsigned((+wire162[(2'h3):(1'h0)]))));
            end
          reg193 = (~reg173);
          reg194 = reg182;
          reg195 <= $unsigned($signed($unsigned(((reg184 ?
              reg179 : forvar189) & $signed(wire162)))));
          for (forvar196 = (1'h0); (forvar196 < (2'h2)); forvar196 = (forvar196 + (1'h1)))
            begin
              reg197 <= reg170[(1'h0):(1'h0)];
              reg198 <= reg170;
              reg199 <= ((&((&{reg179, (8'hba)}) << reg178)) ?
                  reg180[(2'h2):(2'h2)] : wire165[(1'h1):(1'h1)]);
              reg200 <= reg193[(4'hd):(3'h5)];
            end
        end
    end
  always
    @(posedge clk) begin
      reg201 <= (($unsigned((|reg198)) ?
              ({reg187} << $signed((forvar177 <<< reg175))) : reg173) ?
          $signed($signed((((7'h41) && forvar189) ?
              (^reg194) : reg178[(3'h5):(1'h1)]))) : forvar196);
    end
  assign wire202 = (~|reg192[(1'h0):(1'h0)]);
  assign wire203 = forvar189;
  always
    @(posedge clk) begin
      reg204 = $signed(wire161[(4'hf):(3'h4)]);
      reg205 <= ((wire162[(3'h4):(3'h4)] ?
          $unsigned($signed(wire165)) : (8'hbf)) ^~ $signed((($unsigned(reg200) ^ (wire162 << reg178)) >> ((wire164 <= (8'ha0)) >>> (reg185 * wire172)))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module31
#( parameter param156 = {(^~{(&(|(8'ha1))), ({(7'h44), (8'ha7)} ? ((7'h42) ? (8'hae) : (8'hbf)) : (^(8'ha1)))})} )
(y, clk, wire35, wire34, wire33, wire32);
  output wire [(32'h2c5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h9):(1'h0)] wire35;
  input wire signed [(3'h5):(1'h0)] wire34;
  input wire [(4'hc):(1'h0)] wire33;
  input wire [(5'h12):(1'h0)] wire32;
  reg signed [(4'hb):(1'h0)] reg155 = (1'h0);
  reg [(5'h11):(1'h0)] reg154 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg153 = (1'h0);
  reg signed [(4'he):(1'h0)] reg152 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg151 = (1'h0);
  reg [(4'hf):(1'h0)] forvar150 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg149 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg148 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg147 = (1'h0);
  reg [(3'h6):(1'h0)] reg146 = (1'h0);
  reg [(4'hd):(1'h0)] reg145 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire144;
  wire [(4'hb):(1'h0)] wire142;
  wire signed [(4'h8):(1'h0)] wire80;
  reg signed [(4'hd):(1'h0)] reg79 = (1'h0);
  reg [(4'hd):(1'h0)] reg78 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg77 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg76 = (1'h0);
  reg [(5'h15):(1'h0)] reg75 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg74 = (1'h0);
  reg [(3'h4):(1'h0)] forvar73 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire72;
  wire signed [(5'h15):(1'h0)] wire71;
  wire signed [(4'hc):(1'h0)] wire70;
  reg signed [(4'hc):(1'h0)] reg69 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar68 = (1'h0);
  reg [(5'h10):(1'h0)] reg67 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg66 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg65 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg64 = (1'h0);
  reg [(3'h6):(1'h0)] reg63 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg62 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar61 = (1'h0);
  reg [(4'he):(1'h0)] reg60 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar59 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg58 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg57 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire56;
  reg signed [(5'h10):(1'h0)] reg55 = (1'h0);
  reg [(5'h15):(1'h0)] reg54 = (1'h0);
  reg [(5'h10):(1'h0)] reg53 = (1'h0);
  reg [(4'hc):(1'h0)] reg52 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar51 = (1'h0);
  wire [(4'h9):(1'h0)] wire50;
  reg signed [(4'h8):(1'h0)] reg49 = (1'h0);
  reg [(4'hd):(1'h0)] reg48 = (1'h0);
  reg [(3'h7):(1'h0)] reg47 = (1'h0);
  reg signed [(4'he):(1'h0)] reg46 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg45 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg44 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar43 = (1'h0);
  reg [(3'h5):(1'h0)] reg42 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg41 = (1'h0);
  reg [(5'h14):(1'h0)] reg40 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg39 = (1'h0);
  wire [(4'hd):(1'h0)] wire38;
  reg [(3'h6):(1'h0)] reg37 = (1'h0);
  reg [(3'h6):(1'h0)] reg36 = (1'h0);
  assign y = {reg155,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 forvar150,
                 reg149,
                 reg148,
                 reg147,
                 reg146,
                 reg145,
                 wire144,
                 wire142,
                 wire80,
                 reg79,
                 reg78,
                 reg77,
                 reg76,
                 reg75,
                 reg74,
                 forvar73,
                 wire72,
                 wire71,
                 wire70,
                 reg69,
                 forvar68,
                 reg67,
                 reg66,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 forvar61,
                 reg60,
                 forvar59,
                 reg58,
                 reg57,
                 wire56,
                 reg55,
                 reg54,
                 reg53,
                 reg52,
                 forvar51,
                 wire50,
                 reg49,
                 reg48,
                 reg47,
                 reg46,
                 reg45,
                 reg44,
                 forvar43,
                 reg42,
                 reg41,
                 reg40,
                 reg39,
                 wire38,
                 reg37,
                 reg36,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg36 <= ((~|wire33) << $signed((($signed(wire32) >> (wire35 ?
              (8'hbc) : wire34)) ?
          $unsigned(wire32[(3'h7):(3'h5)]) : ($unsigned(wire33) ^ $signed(wire33)))));
    end
  always
    @(posedge clk) begin
      reg37 <= (((|(&((8'hbc) <= reg36))) > {($signed(wire35) ^ $signed(reg36))}) * $unsigned({((wire34 & (8'hb5)) | $signed((8'h9c)))}));
    end
  assign wire38 = (8'hbf);
  always
    @(posedge clk) begin
      reg39 <= ($unsigned($unsigned($unsigned($signed(wire32)))) != $signed(reg37));
      reg40 <= wire38[(4'h8):(3'h6)];
    end
  always
    @(posedge clk) begin
      reg41 <= reg40;
      reg42 <= (wire32 | (wire38 ? (+reg41) : {$signed((reg36 <= reg39))}));
      for (forvar43 = (1'h0); (forvar43 < (2'h3)); forvar43 = (forvar43 + (1'h1)))
        begin
          reg44 <= (~&wire32[(5'h10):(4'hc)]);
          reg45 = (|((-$unsigned(wire33)) ?
              $unsigned($unsigned((wire32 ?
                  reg39 : (8'hbc)))) : (wire35[(1'h0):(1'h0)] ^~ wire35[(4'h8):(2'h3)])));
        end
      reg46 <= (~^$signed((7'h42)));
    end
  always
    @(posedge clk) begin
      reg47 <= reg36[(2'h2):(1'h1)];
      reg48 = reg36;
      reg49 <= $signed($signed((~&$unsigned((reg48 + wire32)))));
    end
  assign wire50 = {(reg40 << wire38[(4'hd):(4'h9)])};
  always
    @(posedge clk) begin
      for (forvar51 = (1'h0); (forvar51 < (2'h2)); forvar51 = (forvar51 + (1'h1)))
        begin
          reg52 <= $unsigned(($signed(((!reg47) + (+forvar51))) ?
              (^$signed($unsigned(wire50))) : (^{reg48})));
        end
      reg53 <= {(reg41 < ($signed(((8'ha7) ? reg44 : forvar51)) ?
              reg41 : reg45)),
          reg42};
      reg54 = reg44[(4'h8):(3'h6)];
      reg55 <= ((^~$unsigned(reg36[(2'h3):(2'h3)])) | $unsigned({$signed($signed((8'hb4)))}));
    end
  assign wire56 = ($unsigned(($unsigned(reg49) ?
                      (reg36[(3'h5):(3'h5)] ~^ wire33[(4'h9):(2'h2)]) : reg53[(4'h9):(3'h5)])) <<< (~^$signed((&wire33[(4'h9):(2'h3)]))));
  always
    @(posedge clk) begin
      reg57 <= {$unsigned({(~^$unsigned(reg45))}), wire56[(3'h7):(3'h5)]};
      reg58 <= (reg42 > reg39);
      for (forvar59 = (1'h0); (forvar59 < (2'h2)); forvar59 = (forvar59 + (1'h1)))
        begin
          reg60 <= reg42;
          for (forvar61 = (1'h0); (forvar61 < (3'h4)); forvar61 = (forvar61 + (1'h1)))
            begin
              reg62 <= reg45[(3'h5):(1'h1)];
              reg63 <= ((reg54[(4'ha):(3'h4)] ?
                      reg41[(4'hf):(2'h2)] : (|reg37)) ?
                  {$unsigned({$unsigned(forvar61)})} : ($unsigned($unsigned(reg39)) ?
                      $unsigned((((8'hb9) || wire34) ^~ (forvar61 ?
                          reg48 : reg57))) : $signed(((reg52 + wire50) ?
                          (wire34 ? reg48 : reg39) : $unsigned(reg60)))));
            end
          reg64 = forvar51;
          reg65 <= $signed($unsigned((reg63[(3'h6):(3'h5)] ?
              $unsigned({wire50}) : ({reg55, wire34} ?
                  $unsigned(reg47) : {reg63}))));
          reg66 = reg60[(4'hb):(3'h5)];
        end
      reg67 <= $signed({$signed({reg49[(2'h2):(1'h0)], (reg60 - reg64)}),
          ($unsigned($unsigned(reg66)) >>> ($unsigned(reg66) - (7'h42)))});
    end
  always
    @(posedge clk) begin
      for (forvar68 = (1'h0); (forvar68 < (1'h1)); forvar68 = (forvar68 + (1'h1)))
        begin
          reg69 <= reg36[(2'h3):(2'h3)];
        end
    end
  assign wire70 = $unsigned($unsigned((reg65 || {((8'ha4) & reg49),
                      (wire56 > reg42)})));
  assign wire71 = $signed(reg64);
  assign wire72 = reg48;
  always
    @(posedge clk) begin
      for (forvar73 = (1'h0); (forvar73 < (3'h4)); forvar73 = (forvar73 + (1'h1)))
        begin
          reg74 <= forvar51[(4'hc):(4'ha)];
          reg75 = ((((8'hb1) ?
              forvar43 : reg46[(1'h1):(1'h0)]) <= ($unsigned($unsigned(forvar61)) ^ reg49[(1'h0):(1'h0)])) | $unsigned((($signed(forvar43) ?
              reg39 : ((8'ha0) ? reg48 : reg39)) | (reg40 ?
              $signed(reg52) : (reg63 ? reg47 : reg55)))));
          reg76 <= $signed($signed($unsigned((|$signed(wire34)))));
          reg77 <= (~|reg36);
          reg78 <= reg39[(5'h13):(4'hb)];
        end
      reg79 <= (reg54 ?
          ({reg75, reg66} == ((-{forvar51,
              wire33}) < reg67[(3'h6):(3'h6)])) : $signed(($signed(reg37[(3'h6):(2'h2)]) >>> ((reg64 && reg60) ^~ $unsigned(wire38)))));
    end
  assign wire80 = (^~reg42);
  module81 modinst143 (.wire85(reg67), .clk(clk), .wire83(reg41), .wire82(reg78), .wire84(forvar68), .y(wire142));
  assign wire144 = (~reg53[(4'h8):(3'h6)]);
  always
    @(posedge clk) begin
      reg145 <= $signed(reg52);
      reg146 <= $unsigned((($unsigned((!reg39)) ?
              $signed(reg36) : $unsigned(reg145[(4'hc):(3'h4)])) ?
          $signed((^~{reg49})) : $signed((~^{reg145}))));
      reg147 = (((^(wire80[(4'h8):(3'h7)] ?
              forvar51[(3'h6):(3'h4)] : $unsigned((8'had)))) >>> ((8'ha2) ?
              $unsigned((8'h9f)) : $unsigned((~wire38)))) ?
          reg54 : reg78[(2'h2):(1'h1)]);
      reg148 <= $signed($unsigned((8'hb2)));
    end
  always
    @(posedge clk) begin
      reg149 = (!{reg39[(4'ha):(3'h5)]});
      for (forvar150 = (1'h0); (forvar150 < (2'h3)); forvar150 = (forvar150 + (1'h1)))
        begin
          reg151 = forvar73;
          reg152 <= reg149[(2'h3):(1'h1)];
          reg153 <= wire56[(1'h0):(1'h0)];
          reg154 <= $unsigned((8'h9d));
        end
      reg155 <= ((reg39[(4'hf):(4'h8)] ?
              {((8'hb6) ? $unsigned(reg154) : (~|(8'hba)))} : reg52) ?
          $signed($unsigned(reg36[(1'h1):(1'h1)])) : $signed({reg153}));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module81
#( parameter param140 = ({((((8'had) < (8'hac)) * (!(7'h44))) ? {((8'hb1) <<< (8'ha6))} : {((8'hb5) ? (7'h40) : (8'hb2))})} ? (((((8'hb7) ? (8'hb2) : (8'h9d)) > ((8'hae) ? (8'hb7) : (8'hb5))) ? (((7'h44) || (8'ha5)) || ((7'h41) ? (8'hbf) : (8'hb5))) : {((8'hbe) ? (8'hb6) : (7'h44)), (^~(8'hb9))}) ? {({(8'ha2)} ? ((8'hb1) ? (8'hbb) : (8'haf)) : (~(8'ha8))), ((+(8'ha7)) + ((8'hb2) ~^ (8'h9e)))} : ((^~{(8'ha0), (8'ha4)}) ? (8'hba) : (~^((8'haa) ^ (8'ha8))))) : ((&(((8'ha2) != (7'h40)) ? {(8'ha7)} : ((8'hb5) && (8'hbe)))) & (^{((7'h41) ? (7'h40) : (8'hae)), {(8'hb2), (8'hb0)}})))
, parameter param141 = (^(((7'h42) >> (-(-param140))) || (param140 >>> (param140 >= (~|param140))))) )
(y, clk, wire85, wire84, wire83, wire82);
  output wire [(32'h25c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire85;
  input wire signed [(2'h3):(1'h0)] wire84;
  input wire [(2'h3):(1'h0)] wire83;
  input wire [(4'hb):(1'h0)] wire82;
  wire [(4'hb):(1'h0)] wire139;
  wire signed [(4'hf):(1'h0)] wire138;
  reg signed [(3'h6):(1'h0)] reg137 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg136 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg135 = (1'h0);
  reg [(2'h2):(1'h0)] reg134 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg133 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg132 = (1'h0);
  reg [(5'h13):(1'h0)] reg131 = (1'h0);
  reg [(5'h11):(1'h0)] forvar130 = (1'h0);
  reg [(2'h2):(1'h0)] reg129 = (1'h0);
  reg [(4'hc):(1'h0)] reg128 = (1'h0);
  reg [(3'h4):(1'h0)] reg127 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg126 = (1'h0);
  reg [(5'h15):(1'h0)] reg125 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg124 = (1'h0);
  reg [(2'h2):(1'h0)] reg123 = (1'h0);
  reg [(5'h14):(1'h0)] reg122 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar121 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg120 = (1'h0);
  reg [(4'hc):(1'h0)] reg119 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg118 = (1'h0);
  reg [(4'hd):(1'h0)] reg117 = (1'h0);
  reg [(4'hd):(1'h0)] reg116 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg115 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg114 = (1'h0);
  reg [(4'hc):(1'h0)] forvar113 = (1'h0);
  reg [(3'h4):(1'h0)] reg112 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg111 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire110;
  reg signed [(5'h13):(1'h0)] reg109 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg108 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg107 = (1'h0);
  reg [(4'hb):(1'h0)] reg106 = (1'h0);
  wire [(5'h15):(1'h0)] wire105;
  wire signed [(3'h4):(1'h0)] wire104;
  wire [(5'h12):(1'h0)] wire103;
  wire signed [(4'ha):(1'h0)] wire102;
  reg signed [(2'h3):(1'h0)] reg101 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar100 = (1'h0);
  reg [(4'h8):(1'h0)] reg99 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg98 = (1'h0);
  reg [(4'hb):(1'h0)] reg97 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg96 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg95 = (1'h0);
  reg [(5'h12):(1'h0)] reg94 = (1'h0);
  reg [(5'h15):(1'h0)] reg93 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar92 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg91 = (1'h0);
  reg [(3'h6):(1'h0)] forvar90 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg89 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg88 = (1'h0);
  reg [(3'h4):(1'h0)] reg87 = (1'h0);
  wire [(5'h11):(1'h0)] wire86;
  assign y = {wire139,
                 wire138,
                 reg137,
                 reg136,
                 reg135,
                 reg134,
                 reg133,
                 reg132,
                 reg131,
                 forvar130,
                 reg129,
                 reg128,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 forvar121,
                 reg120,
                 reg119,
                 reg118,
                 reg117,
                 reg116,
                 reg115,
                 reg114,
                 forvar113,
                 reg112,
                 reg111,
                 wire110,
                 reg109,
                 reg108,
                 reg107,
                 reg106,
                 wire105,
                 wire104,
                 wire103,
                 wire102,
                 reg101,
                 forvar100,
                 reg99,
                 reg98,
                 reg97,
                 reg96,
                 reg95,
                 reg94,
                 reg93,
                 forvar92,
                 reg91,
                 forvar90,
                 reg89,
                 reg88,
                 reg87,
                 wire86,
                 (1'h0)};
  assign wire86 = $signed($unsigned({(~|(~|wire83)), {(wire82 | wire85)}}));
  always
    @(posedge clk) begin
      reg87 <= wire86[(2'h3):(2'h3)];
      reg88 = $unsigned((~^$signed((&wire83))));
      reg89 = wire84;
      for (forvar90 = (1'h0); (forvar90 < (1'h0)); forvar90 = (forvar90 + (1'h1)))
        begin
          reg91 <= wire82[(1'h0):(1'h0)];
          for (forvar92 = (1'h0); (forvar92 < (2'h2)); forvar92 = (forvar92 + (1'h1)))
            begin
              reg93 <= (({$unsigned((wire82 ? (8'ha6) : wire82))} ?
                  (+((reg87 * wire82) ?
                      {wire86,
                          (8'hb2)} : $unsigned((8'haf)))) : reg88) ~^ wire84);
              reg94 = wire86[(4'hb):(4'h9)];
              reg95 = reg93;
              reg96 <= wire85[(1'h1):(1'h0)];
            end
          reg97 <= {(($unsigned((~|(8'haf))) * (~|$unsigned((8'hbd)))) != (+reg87))};
          reg98 <= forvar90[(3'h6):(3'h5)];
        end
      reg99 <= (($unsigned($signed((-wire86))) ?
          {$unsigned(wire83)} : reg94) < {(+$unsigned($unsigned(reg89))),
          reg95[(4'h9):(1'h0)]});
    end
  always
    @(posedge clk) begin
      for (forvar100 = (1'h0); (forvar100 < (2'h3)); forvar100 = (forvar100 + (1'h1)))
        begin
          reg101 <= forvar100[(3'h4):(1'h1)];
        end
    end
  assign wire102 = ((($unsigned((reg95 < (8'ha1))) && ($signed((8'hbc)) ?
                           (wire85 >>> (8'ha5)) : reg87[(3'h4):(3'h4)])) <<< ((^~(reg97 ?
                               reg89 : (8'hbc))) ?
                           ({(8'hac), reg96} ?
                               $unsigned(wire84) : (~&wire85)) : $signed(reg88[(1'h0):(1'h0)]))) ?
                       {forvar92[(2'h2):(1'h1)]} : (8'hb8));
  assign wire103 = $unsigned($signed((8'ha6)));
  assign wire104 = reg91[(2'h3):(1'h1)];
  assign wire105 = ((((8'ha9) ?
                           ({wire102, reg91} ?
                               $unsigned(reg93) : (reg87 != forvar90)) : {(~|reg96)}) ?
                       reg95[(4'h9):(1'h0)] : ({{forvar92}} | wire82)) ~^ (^$unsigned(reg93)));
  always
    @(posedge clk) begin
      reg106 <= reg91;
      reg107 <= ((reg94[(3'h4):(2'h3)] ?
              $signed($unsigned((reg94 ?
                  forvar90 : reg99))) : $signed(($unsigned(reg94) ?
                  $unsigned(reg94) : (wire105 ? (8'hbf) : reg91)))) ?
          $signed($signed(reg89[(2'h3):(1'h1)])) : (&$unsigned(reg94[(4'he):(4'h9)])));
      reg108 <= $unsigned({$unsigned(wire102),
          (^~($signed(reg95) | $unsigned(forvar100)))});
      reg109 <= (reg108 ? $signed((8'hb9)) : reg89[(1'h1):(1'h0)]);
    end
  assign wire110 = {({{$signed(reg94)},
                           $signed($unsigned(reg93))} >> {wire83})};
  always
    @(posedge clk) begin
      reg111 <= $signed((&$unsigned(reg94)));
    end
  always
    @(posedge clk) begin
      reg112 = $unsigned($unsigned($unsigned($signed(reg91))));
      for (forvar113 = (1'h0); (forvar113 < (2'h2)); forvar113 = (forvar113 + (1'h1)))
        begin
          reg114 <= ($signed(reg97[(4'h9):(2'h2)]) ?
              (~&(8'hbe)) : $unsigned(reg96[(4'h9):(1'h0)]));
          reg115 <= (~&(8'ha4));
          reg116 = ($unsigned((($unsigned(reg94) ?
              (reg101 ? (8'ha6) : (8'ha9)) : reg107) * reg89)) > (8'h9d));
          reg117 <= $unsigned(reg97[(4'ha):(3'h6)]);
          reg118 <= (~reg94);
        end
      reg119 = ((&reg107[(3'h6):(2'h3)]) || $signed((8'hab)));
      reg120 <= wire83[(1'h0):(1'h0)];
    end
  always
    @(posedge clk) begin
      for (forvar121 = (1'h0); (forvar121 < (3'h4)); forvar121 = (forvar121 + (1'h1)))
        begin
          reg122 <= (~|(($unsigned((reg88 ? reg117 : reg107)) ?
              $signed({forvar92}) : reg99) || $signed(reg119)));
          reg123 <= reg118;
          reg124 <= (({((reg112 || reg99) ? reg99 : wire102[(1'h0):(1'h0)]),
                      ($signed((8'hb9)) ? (8'hb9) : $unsigned(reg114))} ?
                  (&{wire104[(2'h3):(1'h1)], (^reg115)}) : (wire103 ?
                      reg106[(4'h9):(1'h0)] : $unsigned($unsigned(reg91)))) ?
              (8'ha7) : (reg89[(3'h4):(3'h4)] ?
                  $signed((8'hb9)) : $signed(wire86)));
        end
      reg125 = $unsigned((+wire86));
      reg126 <= reg124[(2'h3):(2'h3)];
      reg127 <= reg115[(1'h0):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg128 <= wire103[(4'hb):(2'h2)];
      reg129 <= $signed($signed(((((8'hb2) ? forvar113 : wire104) ?
              $signed(wire82) : wire105) ?
          (~^wire85) : (~^forvar100))));
      for (forvar130 = (1'h0); (forvar130 < (3'h4)); forvar130 = (forvar130 + (1'h1)))
        begin
          reg131 <= reg119[(4'h8):(3'h5)];
          reg132 <= $signed(($unsigned($unsigned((wire86 ?
                  reg112 : forvar113))) ?
              forvar90[(3'h6):(3'h5)] : $signed(reg89)));
          reg133 <= ($unsigned(({(reg126 ?
                  (7'h40) : (8'h9e))} * reg98)) << wire82[(1'h0):(1'h0)]);
          if ((^~(~^(8'ha2))))
            begin
              reg134 = ((~|$signed($unsigned((~(7'h44))))) - (reg107[(2'h2):(2'h2)] != ((^((8'ha4) != reg115)) < reg89)));
            end
          else
            begin
              reg134 <= $signed(forvar90);
              reg135 <= $signed({$unsigned((reg101 ?
                      $unsigned(reg87) : $unsigned(reg89)))});
            end
          reg136 <= $signed(((7'h41) != $signed(reg98[(3'h7):(3'h6)])));
        end
      reg137 = $signed((-wire102[(2'h3):(1'h0)]));
    end
  assign wire138 = forvar100[(2'h2):(1'h0)];
  assign wire139 = (~|reg111);
endmodule