(* use_dsp48="no" *) (* use_dsp="no" *) module top
#( parameter param1476 = ((+{(((8'hb5) ? (8'ha4) : (8'hb9)) ^ (~^(8'hb0)))}) ? ((|{(~^(8'hb0)), ((8'hb8) | (8'hb1))}) ? (((~|(8'hb5)) | ((8'hb0) || (8'ha7))) ? (^~((7'h43) & (8'hab))) : ((8'h9c) ? ((8'hbf) ? (8'hae) : (8'ha4)) : ((7'h44) << (8'hb1)))) : ((!(~^(8'h9f))) ? (~((8'hae) ? (8'hb4) : (8'ha9))) : ((+(8'h9e)) ? (-(8'ha6)) : ((8'ha0) ? (8'hae) : (8'haa))))) : ((|{(|(8'hbb)), ((8'hb5) ? (8'hbc) : (8'hb9))}) != (&(((8'hb4) ? (8'ha4) : (7'h41)) ? ((8'ha5) ? (8'ha8) : (8'hbb)) : (!(7'h42))))))
, parameter param1477 = {(|param1476)} )
(y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h1cb):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h9):(1'h0)] wire3;
  input wire [(3'h4):(1'h0)] wire2;
  input wire signed [(5'h11):(1'h0)] wire1;
  input wire signed [(2'h2):(1'h0)] wire0;
  wire signed [(5'h14):(1'h0)] wire1447;
  wire signed [(3'h6):(1'h0)] wire15;
  wire signed [(5'h13):(1'h0)] wire14;
  wire [(4'hd):(1'h0)] wire13;
  wire [(5'h15):(1'h0)] wire12;
  wire [(3'h4):(1'h0)] wire11;
  reg signed [(3'h6):(1'h0)] reg10 = (1'h0);
  reg [(5'h12):(1'h0)] reg9 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg8 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar7 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6 = (1'h0);
  reg [(4'he):(1'h0)] reg5 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4 = (1'h0);
  reg [(4'h9):(1'h0)] reg1449 = (1'h0);
  reg [(3'h4):(1'h0)] reg1450 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1451 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire1452;
  wire signed [(4'hc):(1'h0)] wire1453;
  wire [(2'h3):(1'h0)] wire1454;
  wire signed [(3'h7):(1'h0)] wire1455;
  reg signed [(5'h14):(1'h0)] reg1456 = (1'h0);
  reg [(5'h15):(1'h0)] reg1457 = (1'h0);
  reg [(3'h7):(1'h0)] reg1458 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire1459;
  reg [(5'h12):(1'h0)] reg1460 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1461 = (1'h0);
  reg [(4'h9):(1'h0)] reg1462 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1463 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1464 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1465 = (1'h0);
  reg [(4'hf):(1'h0)] reg1466 = (1'h0);
  reg [(2'h3):(1'h0)] reg1467 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1468 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1469 = (1'h0);
  reg [(5'h14):(1'h0)] reg1470 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1471 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1472 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire1473;
  wire [(4'hd):(1'h0)] wire1474;
  assign y = {wire1447,
                 wire15,
                 wire14,
                 wire13,
                 wire12,
                 wire11,
                 reg10,
                 reg9,
                 reg8,
                 forvar7,
                 reg6,
                 reg5,
                 reg4,
                 reg1449,
                 reg1450,
                 reg1451,
                 wire1452,
                 wire1453,
                 wire1454,
                 wire1455,
                 reg1456,
                 reg1457,
                 reg1458,
                 wire1459,
                 reg1460,
                 reg1461,
                 reg1462,
                 forvar1463,
                 reg1464,
                 reg1465,
                 reg1466,
                 reg1467,
                 forvar1468,
                 reg1469,
                 reg1470,
                 reg1471,
                 reg1472,
                 wire1473,
                 wire1474,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg4 = $signed(($unsigned($signed(wire3[(1'h0):(1'h0)])) <<< wire0[(1'h1):(1'h1)]));
      reg5 <= $signed((wire3[(2'h2):(1'h0)] ~^ {{$signed((8'hb3))}}));
      reg6 <= ((wire0[(2'h2):(1'h0)] ?
          reg4 : $unsigned((~(reg5 && wire2)))) || $unsigned((~&(wire0 ?
          wire2 : (wire0 ? reg4 : (8'hac))))));
      for (forvar7 = (1'h0); (forvar7 < (1'h1)); forvar7 = (forvar7 + (1'h1)))
        begin
          reg8 <= $unsigned(reg6);
          reg9 <= (8'ha0);
          reg10 = ((forvar7 ^~ ((+wire3[(2'h3):(1'h0)]) & {(wire3 ^ reg9)})) == (^~$unsigned($signed(reg8[(3'h5):(1'h1)]))));
        end
    end
  assign wire11 = wire0;
  assign wire12 = $signed((&$unsigned({(wire0 - wire0), $unsigned((8'hbd))})));
  assign wire13 = wire11[(1'h1):(1'h1)];
  assign wire14 = $signed((~((-$unsigned(wire2)) ?
                      ($signed(wire0) * $signed(reg4)) : $unsigned($unsigned(wire0)))));
  assign wire15 = (wire2 | wire13[(1'h1):(1'h1)]);
  module16 modinst1448 (.clk(clk), .wire19(reg9), .wire18(wire13), .wire20(wire3), .wire21(reg4), .wire17(forvar7), .y(wire1447));
  always
    @(posedge clk) begin
      reg1449 <= $signed(wire2[(2'h3):(2'h2)]);
      reg1450 <= $signed({$signed((+wire15)), reg1449});
      reg1451 <= $signed(((wire0 <= {forvar7[(1'h0):(1'h0)]}) ?
          $unsigned((~$unsigned(reg1450))) : (($unsigned(reg1449) >> $unsigned((8'ha5))) > $signed($unsigned(wire1447)))));
    end
  assign wire1452 = wire11;
  assign wire1453 = (forvar7 ? wire15[(1'h1):(1'h0)] : reg8);
  assign wire1454 = $signed($unsigned(reg8));
  assign wire1455 = (~^{$signed($signed($signed(wire0)))});
  always
    @(posedge clk) begin
      reg1456 <= {($signed((wire1[(4'hd):(4'hd)] ?
              $unsigned(wire14) : ((8'h9e) << wire1))) < $unsigned($signed((-wire3))))};
      reg1457 <= reg5[(1'h1):(1'h0)];
      reg1458 <= wire1453[(4'h8):(3'h7)];
    end
  assign wire1459 = $signed($unsigned(((8'ha6) - (+{reg6}))));
  always
    @(posedge clk) begin
      reg1460 <= (&wire11);
      reg1461 <= $signed($signed({{(wire15 ? wire1453 : wire2)}}));
      reg1462 <= $unsigned($unsigned(wire14));
      for (forvar1463 = (1'h0); (forvar1463 < (1'h0)); forvar1463 = (forvar1463 + (1'h1)))
        begin
          reg1464 <= ($unsigned((wire13[(2'h2):(1'h1)] ?
              ($unsigned(forvar1463) != (wire1453 ?
                  wire1 : reg8)) : (reg8 != reg1451[(2'h3):(2'h2)]))) || forvar7[(2'h3):(2'h3)]);
          reg1465 = ((~&(reg1450[(2'h2):(1'h1)] ?
              ((&reg1450) ?
                  {(8'hb4)} : reg1449) : wire1459[(3'h5):(1'h1)])) >> (($signed((reg6 ?
                      forvar7 : wire1453)) ?
                  reg1456 : $signed((reg1450 <<< reg1449))) ?
              (~|((reg5 <<< reg1462) ?
                  (reg1462 || wire2) : (reg1450 ?
                      reg4 : wire13))) : $signed($signed($unsigned(wire3)))));
          reg1466 = $unsigned($unsigned((((forvar7 >> wire13) >= wire1459) != wire1459[(2'h3):(1'h1)])));
          reg1467 <= (~|(wire1452 >= (wire15 * $signed((reg1450 >>> reg1464)))));
          for (forvar1468 = (1'h0); (forvar1468 < (3'h4)); forvar1468 = (forvar1468 + (1'h1)))
            begin
              reg1469 = $unsigned((|wire3[(1'h0):(1'h0)]));
              reg1470 = ($unsigned($signed((((8'ha6) || (8'h9c)) > (wire1452 ?
                      reg1462 : (8'h9f))))) ?
                  (8'hb1) : reg1450);
              reg1471 = {((forvar1468 >>> $unsigned(reg1451)) ?
                      $unsigned((~wire1459[(1'h1):(1'h0)])) : $unsigned((~|wire1453[(3'h4):(3'h4)]))),
                  wire3[(1'h1):(1'h1)]};
              reg1472 = $signed($unsigned(wire11[(3'h4):(2'h3)]));
            end
        end
    end
  assign wire1473 = ((wire3[(2'h2):(1'h1)] ?
                            wire1452[(4'ha):(3'h5)] : wire1452) ?
                        $unsigned($unsigned(({reg1456, reg1456} ^~ (reg1467 ?
                            (8'hb4) : reg1464)))) : reg1465);
  module688 modinst1475 (.wire692(reg1470), .wire693(wire1452), .wire691(reg1471), .clk(clk), .wire689(reg1464), .y(wire1474), .wire690(wire1));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module16
#( parameter param1445 = ((~|{({(8'ha9), (8'hb5)} ? ((8'ha7) ? (8'ha9) : (7'h40)) : {(8'hb8)})}) <<< (8'hbc))
, parameter param1446 = (param1445 > param1445) )
(y, clk, wire21, wire20, wire19, wire18, wire17);
  output wire [(32'h21e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h7):(1'h0)] wire21;
  input wire signed [(4'h9):(1'h0)] wire20;
  input wire [(5'h12):(1'h0)] wire19;
  input wire signed [(4'hd):(1'h0)] wire18;
  input wire signed [(2'h2):(1'h0)] wire17;
  reg [(3'h4):(1'h0)] reg1444 = (1'h0);
  reg [(3'h4):(1'h0)] reg1443 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1442 = (1'h0);
  reg [(3'h6):(1'h0)] reg1433 = (1'h0);
  reg [(5'h14):(1'h0)] reg1441 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1440 = (1'h0);
  reg [(5'h14):(1'h0)] reg1439 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1438 = (1'h0);
  reg [(3'h6):(1'h0)] reg1437 = (1'h0);
  reg [(5'h13):(1'h0)] reg1436 = (1'h0);
  reg [(5'h12):(1'h0)] reg1435 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1434 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1433 = (1'h0);
  reg [(3'h5):(1'h0)] reg1432 = (1'h0);
  wire [(5'h15):(1'h0)] wire1431;
  wire signed [(5'h11):(1'h0)] wire1430;
  wire [(2'h3):(1'h0)] wire1429;
  reg signed [(3'h7):(1'h0)] reg1428 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1427 = (1'h0);
  reg [(4'hd):(1'h0)] reg1426 = (1'h0);
  reg [(4'hb):(1'h0)] reg1425 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1424 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1423 = (1'h0);
  reg [(4'hd):(1'h0)] reg1422 = (1'h0);
  reg [(5'h10):(1'h0)] reg1421 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1420 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire1418;
  wire [(4'hd):(1'h0)] wire794;
  wire signed [(4'h9):(1'h0)] wire793;
  reg [(4'hb):(1'h0)] reg792 = (1'h0);
  reg [(5'h15):(1'h0)] reg791 = (1'h0);
  reg [(4'hd):(1'h0)] reg790 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire789;
  wire signed [(5'h13):(1'h0)] wire787;
  reg signed [(5'h12):(1'h0)] reg34 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg33 = (1'h0);
  reg [(5'h12):(1'h0)] reg32 = (1'h0);
  reg [(4'h9):(1'h0)] reg31 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg30 = (1'h0);
  reg [(5'h12):(1'h0)] reg29 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg28 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg27 = (1'h0);
  reg [(4'ha):(1'h0)] reg26 = (1'h0);
  reg [(3'h7):(1'h0)] reg25 = (1'h0);
  reg [(5'h13):(1'h0)] reg24 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg23 = (1'h0);
  reg [(3'h4):(1'h0)] reg22 = (1'h0);
  assign y = {reg1444,
                 reg1443,
                 reg1442,
                 reg1433,
                 reg1441,
                 reg1440,
                 reg1439,
                 reg1438,
                 reg1437,
                 reg1436,
                 reg1435,
                 reg1434,
                 forvar1433,
                 reg1432,
                 wire1431,
                 wire1430,
                 wire1429,
                 reg1428,
                 reg1427,
                 reg1426,
                 reg1425,
                 reg1424,
                 reg1423,
                 reg1422,
                 reg1421,
                 reg1420,
                 wire1418,
                 wire794,
                 wire793,
                 reg792,
                 reg791,
                 reg790,
                 wire789,
                 wire787,
                 reg34,
                 reg33,
                 reg32,
                 reg31,
                 reg30,
                 reg29,
                 reg28,
                 reg27,
                 reg26,
                 reg25,
                 reg24,
                 reg23,
                 reg22,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg22 <= $signed(({wire20[(1'h0):(1'h0)],
          wire19} - ((wire17[(1'h0):(1'h0)] ?
              (wire20 <<< wire19) : (wire18 ? wire21 : wire19)) ?
          $unsigned($unsigned(wire19)) : (wire18 ?
              ((8'ha1) ? wire20 : (8'ha4)) : (8'h9d)))));
      reg23 <= {{(wire20[(3'h7):(3'h4)] <<< (8'hbe)), reg22},
          ((~(~&$unsigned(wire17))) ?
              (((wire21 ? (7'h41) : wire21) ^~ wire21[(2'h3):(1'h1)]) ?
                  $signed($unsigned(wire19)) : wire18) : reg22)};
      if ((wire20[(3'h6):(2'h2)] ?
          (8'hbf) : ((|(~|reg23)) ?
              ($signed((~&wire20)) >> $signed($unsigned(reg23))) : (reg23 + ($unsigned(wire19) ^ $unsigned(reg22))))))
        begin
          if ($signed(wire21[(2'h2):(1'h1)]))
            begin
              reg24 <= $signed(reg23[(3'h6):(2'h2)]);
              reg25 = {($unsigned($unsigned(((8'hb0) | reg24))) > $signed(wire17)),
                  reg23};
              reg26 <= ((-$signed((~(wire17 ? wire21 : wire18)))) ?
                  wire20 : (8'hbf));
              reg27 <= (((~|(reg26[(4'h9):(3'h5)] * (reg24 ~^ reg23))) ?
                      $signed(((+(8'ha7)) <<< reg22[(1'h1):(1'h0)])) : ($unsigned((wire21 * wire18)) < {$signed(reg23),
                          reg23})) ?
                  $signed(reg26[(2'h3):(2'h2)]) : reg24[(2'h2):(1'h1)]);
              reg28 <= (~|(reg23[(1'h0):(1'h0)] ?
                  (wire17[(1'h0):(1'h0)] < $signed({reg24,
                      wire19})) : (^~$signed((~|reg27)))));
            end
          else
            begin
              reg24 <= $signed(($signed($unsigned(wire17)) | {{reg25, reg23},
                  ((+wire21) - reg25[(2'h3):(1'h1)])}));
              reg25 <= $unsigned(((~|(-$unsigned((8'hb1)))) < $signed($unsigned($signed(reg28)))));
              reg26 <= reg25[(1'h0):(1'h0)];
              reg27 <= (((~^$signed({(7'h40)})) ?
                  (reg27 <= ((8'hb6) & $signed(wire18))) : ($signed({reg27,
                          (8'hb9)}) ?
                      $unsigned(reg28) : (reg24 <= wire17))) && (!$signed((8'ha3))));
            end
          reg29 <= ((8'ha1) ?
              (^~(~^((wire20 ? wire18 : reg26) ?
                  reg27[(1'h1):(1'h0)] : $unsigned(wire18)))) : reg27);
          reg30 <= $unsigned($unsigned((reg22 && ($signed(reg26) ?
              $signed((8'haf)) : wire20))));
          reg31 = (((reg24[(4'ha):(3'h4)] ~^ (reg26[(3'h4):(2'h2)] ?
                      $unsigned(reg24) : reg24[(2'h3):(1'h0)])) ?
                  reg30 : ({wire20,
                      (reg28 ? wire20 : wire17)} + (reg24[(3'h4):(2'h2)] ?
                      wire20[(1'h1):(1'h0)] : wire21[(1'h1):(1'h1)]))) ?
              (((reg24 != (reg25 ? wire17 : reg24)) >> reg27[(4'h9):(2'h2)]) ?
                  reg26[(2'h2):(1'h1)] : (8'ha4)) : $unsigned(wire18[(1'h1):(1'h1)]));
          reg32 = wire21[(3'h6):(3'h5)];
        end
      else
        begin
          reg24 = wire19;
          reg25 = $signed($unsigned(reg22[(2'h2):(1'h0)]));
        end
      reg33 <= $unsigned($signed((8'hb1)));
      reg34 <= wire19;
    end
  module35 modinst788 (.wire37(reg30), .clk(clk), .wire39(reg34), .y(wire787), .wire36(reg24), .wire38(wire18));
  assign wire789 = $signed((wire17 - reg34));
  always
    @(posedge clk) begin
      reg790 <= ((reg30 ?
              $signed(($unsigned(reg25) ?
                  (reg22 == wire17) : $unsigned(wire19))) : (((wire19 != reg25) ?
                  reg31 : (-reg27)) != $signed((~|reg22)))) ?
          ((~wire18[(3'h4):(1'h0)]) < ((wire17[(2'h2):(1'h0)] ?
              $unsigned(wire19) : reg29[(5'h11):(1'h0)]) >> $signed((^~(8'ha4))))) : $unsigned((~(~|{reg24,
              reg30}))));
      reg791 <= ((|reg30[(5'h11):(1'h1)]) < (wire17 << reg30));
      reg792 <= $unsigned(wire17);
    end
  assign wire793 = (($unsigned({$unsigned(reg33),
                           $signed(reg22)}) | $signed($signed($unsigned(reg26)))) ?
                       ($signed(reg30[(3'h7):(2'h2)]) ?
                           reg790 : (~&reg791)) : wire21);
  assign wire794 = $signed(reg791[(4'he):(4'hd)]);
  module795 modinst1419 (.wire799(reg791), .y(wire1418), .wire796(wire19), .wire797(reg30), .clk(clk), .wire798(wire787));
  always
    @(posedge clk) begin
      reg1420 <= ((!(reg791[(5'h14):(4'h8)] ~^ reg790)) < (wire17 ?
          reg25 : ({(~^reg32)} ^ $signed((wire789 ? reg32 : wire789)))));
      reg1421 <= (~&$unsigned(({wire18} ?
          ($signed(reg24) ~^ reg1420) : reg32[(4'hf):(4'hd)])));
      reg1422 = reg29;
    end
  always
    @(posedge clk) begin
      reg1423 = (~|($unsigned(((wire1418 ? reg791 : (7'h42)) >>> (reg1422 ?
              reg27 : reg29))) ?
          $signed(({wire21} ?
              (~&(8'hb7)) : $unsigned(reg30))) : (((8'had) == reg23) ?
              (~^$unsigned((8'hb1))) : $unsigned({reg33, reg28}))));
      reg1424 = $signed((((7'h41) ?
              ({reg790, reg23} | $unsigned(wire787)) : $unsigned((wire1418 ?
                  reg23 : reg1421))) ?
          (~&$signed((-reg1422))) : ($signed($unsigned(reg28)) >= reg30[(4'hf):(4'h9)])));
      reg1425 <= reg25;
    end
  always
    @(posedge clk) begin
      reg1426 <= $signed($signed((^~wire794[(3'h6):(2'h3)])));
      reg1427 <= wire794[(3'h6):(2'h2)];
      reg1428 <= $signed(reg28);
    end
  assign wire1429 = reg1428;
  assign wire1430 = ($unsigned((~^$signed((reg25 <<< reg1421)))) ?
                        $signed((7'h40)) : ({(+{(8'haa)})} ?
                            $unsigned(wire20) : $unsigned(wire20)));
  assign wire1431 = ($signed((({wire787} ?
                            $unsigned((8'hb1)) : $signed((8'hac))) ?
                        reg1423 : $unsigned((wire1430 << wire793)))) <<< (~{{(^~wire793),
                            $signed(wire19)}}));
  always
    @(posedge clk) begin
      reg1432 = wire793;
      if ($signed(((-$signed($signed(reg1423))) ^ $signed(($signed(wire1418) ?
          $unsigned(wire19) : ((8'haa) ? wire19 : wire19))))))
        begin
          for (forvar1433 = (1'h0); (forvar1433 < (2'h2)); forvar1433 = (forvar1433 + (1'h1)))
            begin
              reg1434 <= $unsigned(($unsigned({(reg1420 >>> wire1418),
                      {reg24}}) ?
                  $unsigned(reg1420) : (~(reg1422[(1'h0):(1'h0)] ?
                      (^~reg790) : (reg31 ^ reg34)))));
              reg1435 <= reg1421[(3'h7):(3'h7)];
              reg1436 <= {(~|(8'hb7)), reg1434[(3'h6):(2'h2)]};
              reg1437 <= ({($unsigned($signed(reg1422)) && ({reg1432} ?
                      $unsigned(wire1431) : $unsigned(reg1423))),
                  wire1418[(3'h7):(1'h1)]} != (reg791 >>> (reg28[(2'h3):(2'h3)] + (reg1428[(2'h2):(2'h2)] > reg792))));
              reg1438 = ($unsigned((((wire789 == wire17) != $signed(wire1429)) >> ((^~reg1434) & (!reg792)))) ?
                  ($unsigned($signed($signed(reg1437))) ?
                      reg1436[(3'h4):(2'h3)] : (~|reg1432)) : (($signed($signed(reg22)) ?
                      $unsigned($unsigned(wire17)) : (((8'ha4) ?
                          wire1418 : reg791) ^~ reg1421[(3'h5):(2'h3)])) != $unsigned((-reg1434[(2'h3):(2'h2)]))));
            end
          reg1439 <= (~|(((((8'hb3) || (8'hb1)) ^ $unsigned(reg1432)) + $unsigned(reg1432[(2'h2):(2'h2)])) ?
              wire793 : wire1430));
          reg1440 <= (~|reg1420);
          reg1441 <= wire17;
        end
      else
        begin
          reg1433 <= (^(reg24 ?
              ($unsigned((&reg1432)) && ((wire793 ? wire18 : reg22) ?
                  ((7'h42) != (8'hb4)) : $signed(wire21))) : ((-reg1439[(3'h6):(1'h1)]) ?
                  reg1426[(1'h1):(1'h1)] : reg790)));
          reg1434 <= $unsigned((&($unsigned($unsigned((7'h40))) ?
              (8'hac) : reg22[(2'h3):(1'h1)])));
        end
      reg1442 <= (+((((forvar1433 << forvar1433) ?
              $unsigned(reg792) : $unsigned(reg790)) ?
          wire1429[(2'h3):(1'h0)] : (^~(^~(8'hb2)))) <<< ((8'hbd) ?
          reg1434 : ($unsigned(reg32) == $unsigned(reg1438)))));
      reg1443 <= reg31[(1'h0):(1'h0)];
      reg1444 <= reg1422;
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module795
#( parameter param1416 = (~^({(((8'hb5) <<< (8'hb4)) ? (~(8'ha0)) : (+(7'h42)))} ? (({(8'h9f)} * (^(8'ha0))) >= (((8'hb5) - (8'hb4)) | ((8'hbe) + (8'hbf)))) : (~^{(&(8'hb1))})))
, parameter param1417 = (((param1416 ? (~^(!param1416)) : ((~|(7'h44)) & param1416)) - (&{(param1416 || param1416)})) ? {(^~((param1416 ? param1416 : param1416) >= param1416))} : (((!(^~param1416)) ? {(param1416 ? param1416 : param1416)} : param1416) ^ (((+param1416) ? param1416 : param1416) << (param1416 >> (param1416 ? param1416 : param1416))))) )
(y, clk, wire799, wire798, wire797, wire796);
  output wire [(32'h3b2):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire799;
  input wire signed [(3'h7):(1'h0)] wire798;
  input wire signed [(4'he):(1'h0)] wire797;
  input wire [(4'ha):(1'h0)] wire796;
  wire [(5'h13):(1'h0)] wire1415;
  reg signed [(2'h3):(1'h0)] reg1414 = (1'h0);
  reg [(5'h13):(1'h0)] reg1413 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1412 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1411 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1410 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1409 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1408 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1407 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1406 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1405 = (1'h0);
  reg [(4'hc):(1'h0)] reg1404 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1403 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1402 = (1'h0);
  wire [(4'hc):(1'h0)] wire1401;
  wire [(5'h11):(1'h0)] wire1400;
  wire [(4'hf):(1'h0)] wire1399;
  reg signed [(4'hc):(1'h0)] reg1398 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1397 = (1'h0);
  reg [(4'h8):(1'h0)] reg1396 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1395 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1394 = (1'h0);
  reg [(2'h2):(1'h0)] reg1393 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1392 = (1'h0);
  reg [(3'h7):(1'h0)] reg1391 = (1'h0);
  reg [(3'h4):(1'h0)] reg1390 = (1'h0);
  reg [(3'h5):(1'h0)] reg1389 = (1'h0);
  reg [(4'hd):(1'h0)] reg1388 = (1'h0);
  reg [(4'h8):(1'h0)] reg1387 = (1'h0);
  reg [(2'h2):(1'h0)] reg1386 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1385 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1384 = (1'h0);
  reg [(5'h13):(1'h0)] reg1383 = (1'h0);
  reg [(4'hb):(1'h0)] reg1382 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1381 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1380 = (1'h0);
  reg [(5'h15):(1'h0)] reg1379 = (1'h0);
  wire [(5'h14):(1'h0)] wire1377;
  wire [(4'he):(1'h0)] wire845;
  reg signed [(2'h2):(1'h0)] reg844 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg843 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg842 = (1'h0);
  reg [(5'h13):(1'h0)] forvar841 = (1'h0);
  reg [(2'h3):(1'h0)] reg840 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg839 = (1'h0);
  reg signed [(4'he):(1'h0)] reg838 = (1'h0);
  reg [(5'h10):(1'h0)] reg837 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg836 = (1'h0);
  reg [(3'h5):(1'h0)] reg835 = (1'h0);
  reg [(5'h13):(1'h0)] forvar834 = (1'h0);
  reg [(3'h4):(1'h0)] reg833 = (1'h0);
  reg [(3'h4):(1'h0)] reg832 = (1'h0);
  reg [(3'h5):(1'h0)] reg831 = (1'h0);
  reg [(5'h13):(1'h0)] reg830 = (1'h0);
  reg [(4'hb):(1'h0)] forvar829 = (1'h0);
  reg [(4'h8):(1'h0)] reg828 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg827 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg826 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg825 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg824 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg823 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar822 = (1'h0);
  reg [(5'h12):(1'h0)] forvar821 = (1'h0);
  reg [(5'h10):(1'h0)] reg820 = (1'h0);
  wire [(4'he):(1'h0)] wire819;
  reg [(5'h11):(1'h0)] reg818 = (1'h0);
  reg [(2'h2):(1'h0)] reg817 = (1'h0);
  reg [(3'h6):(1'h0)] reg816 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg815 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg814 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg813 = (1'h0);
  reg [(4'hc):(1'h0)] forvar812 = (1'h0);
  reg [(4'h8):(1'h0)] reg811 = (1'h0);
  wire [(5'h11):(1'h0)] wire810;
  reg [(4'ha):(1'h0)] reg809 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg808 = (1'h0);
  reg [(5'h14):(1'h0)] reg807 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg806 = (1'h0);
  reg [(4'hd):(1'h0)] reg805 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg804 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar803 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg802 = (1'h0);
  reg [(5'h12):(1'h0)] reg801 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg800 = (1'h0);
  assign y = {wire1415,
                 reg1414,
                 reg1413,
                 reg1412,
                 reg1411,
                 forvar1410,
                 reg1409,
                 reg1408,
                 forvar1407,
                 reg1406,
                 reg1405,
                 reg1404,
                 forvar1403,
                 reg1402,
                 wire1401,
                 wire1400,
                 wire1399,
                 reg1398,
                 reg1397,
                 reg1396,
                 forvar1395,
                 reg1394,
                 reg1393,
                 reg1392,
                 reg1391,
                 reg1390,
                 reg1389,
                 reg1388,
                 reg1387,
                 reg1386,
                 reg1385,
                 reg1384,
                 reg1383,
                 reg1382,
                 forvar1381,
                 forvar1380,
                 reg1379,
                 wire1377,
                 wire845,
                 reg844,
                 reg843,
                 reg842,
                 forvar841,
                 reg840,
                 reg839,
                 reg838,
                 reg837,
                 reg836,
                 reg835,
                 forvar834,
                 reg833,
                 reg832,
                 reg831,
                 reg830,
                 forvar829,
                 reg828,
                 reg827,
                 reg826,
                 reg825,
                 reg824,
                 reg823,
                 forvar822,
                 forvar821,
                 reg820,
                 wire819,
                 reg818,
                 reg817,
                 reg816,
                 reg815,
                 reg814,
                 reg813,
                 forvar812,
                 reg811,
                 wire810,
                 reg809,
                 reg808,
                 reg807,
                 reg806,
                 reg805,
                 reg804,
                 forvar803,
                 reg802,
                 reg801,
                 reg800,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg800 <= (wire798[(3'h5):(1'h1)] && ((($signed(wire797) || (wire799 ?
          wire796 : wire798)) != $unsigned((+wire797))) || (((!(8'ha1)) - (wire797 ?
          wire796 : wire796)) | (+(8'hb9)))));
      reg801 <= (~|wire799);
      reg802 <= {reg800};
      for (forvar803 = (1'h0); (forvar803 < (1'h0)); forvar803 = (forvar803 + (1'h1)))
        begin
          reg804 <= (reg801[(3'h6):(1'h1)] ?
              {wire796[(3'h5):(3'h4)]} : wire799[(4'hf):(4'hb)]);
          reg805 <= wire798;
          reg806 <= forvar803;
          reg807 = $signed(wire799);
          reg808 <= ((|reg807[(1'h1):(1'h1)]) || (~|(-(~|$signed(reg802)))));
        end
      reg809 <= $signed((forvar803[(3'h7):(2'h2)] >= $unsigned(reg806[(4'h8):(3'h7)])));
    end
  assign wire810 = reg801[(3'h6):(2'h2)];
  always
    @(posedge clk) begin
      reg811 = ({$unsigned((!(wire799 <= reg800))), wire797} ?
          reg805[(4'ha):(3'h4)] : $signed({{{reg807}, reg805[(4'hc):(3'h5)]}}));
      for (forvar812 = (1'h0); (forvar812 < (3'h4)); forvar812 = (forvar812 + (1'h1)))
        begin
          reg813 <= wire798[(2'h3):(2'h2)];
          reg814 <= ((^wire810) && wire797);
          reg815 <= $unsigned($unsigned((8'hbe)));
        end
      reg816 = $unsigned($signed((((+(8'h9c)) || (wire798 ? reg800 : wire799)) ?
          reg806[(3'h7):(1'h0)] : reg808[(1'h0):(1'h0)])));
      reg817 <= (reg808[(4'h9):(3'h5)] + ((8'hb6) ?
          $signed(({(8'ha4), reg816} ?
              $unsigned((8'hbb)) : reg807[(4'hb):(3'h5)])) : ((&wire799[(3'h5):(2'h3)]) ?
              reg801[(1'h0):(1'h0)] : wire799)));
      reg818 = wire799;
    end
  assign wire819 = $signed(((&$unsigned((!(8'hb6)))) - $signed($signed((wire799 ^~ forvar803)))));
  always
    @(posedge clk) begin
      reg820 <= $unsigned({(-((wire796 ?
              reg801 : (8'h9e)) + reg804[(3'h5):(2'h3)])),
          $signed(wire799)});
    end
  always
    @(posedge clk) begin
      for (forvar821 = (1'h0); (forvar821 < (1'h0)); forvar821 = (forvar821 + (1'h1)))
        begin
          for (forvar822 = (1'h0); (forvar822 < (2'h2)); forvar822 = (forvar822 + (1'h1)))
            begin
              reg823 <= (^~((((reg807 ^~ wire798) >= (reg813 > reg808)) ?
                      (((7'h44) || forvar812) ?
                          $unsigned(reg809) : reg806[(4'h8):(3'h4)]) : $signed({reg817})) ?
                  (8'ha1) : $unsigned($signed({reg816}))));
              reg824 <= {$signed({((&reg801) != wire798[(3'h5):(1'h0)])})};
              reg825 = ((|$unsigned(((reg800 ? reg813 : (7'h44)) ?
                  $unsigned(forvar822) : ((8'ha0) ^ reg820)))) > ((|((~|reg818) ?
                  $signed(reg815) : (-reg818))) <<< ((~((8'hae) ?
                      reg805 : (8'hb1))) ?
                  (~&$unsigned(reg817)) : (~^$unsigned(reg818)))));
              reg826 <= (!reg809);
            end
          reg827 = {forvar822[(3'h5):(2'h3)],
              (reg813 ~^ $signed($signed((reg809 ? forvar821 : reg826))))};
          reg828 <= (^reg814);
        end
      for (forvar829 = (1'h0); (forvar829 < (3'h4)); forvar829 = (forvar829 + (1'h1)))
        begin
          reg830 <= (-reg805[(4'hb):(1'h0)]);
        end
      reg831 <= wire797;
    end
  always
    @(posedge clk) begin
      reg832 = $signed((~^(reg811 ? forvar822 : (|$signed(reg800)))));
    end
  always
    @(posedge clk) begin
      reg833 <= ((((-(wire796 << reg804)) > ({(8'hae),
                  reg800} <= $signed(reg824))) ?
              (|((|(8'hb2)) <= wire819)) : (reg824 ?
                  reg830 : (~(forvar821 ? forvar822 : reg827)))) ?
          $unsigned(((forvar829 + $signed(reg828)) >> (reg824 ?
              $signed((7'h41)) : (~reg807)))) : (reg815[(4'ha):(1'h0)] ?
              ({$signed(reg830)} ?
                  (reg800 ?
                      (forvar812 ?
                          (7'h44) : wire810) : $unsigned(reg814)) : {(-reg801),
                      $signed(forvar812)}) : (~^((wire819 >= reg817) << (~|(8'hb0))))));
      for (forvar834 = (1'h0); (forvar834 < (3'h4)); forvar834 = (forvar834 + (1'h1)))
        begin
          reg835 <= $signed($unsigned(forvar803));
          reg836 <= $signed((8'hab));
          reg837 = ($unsigned(reg809) << (reg830 * reg818[(1'h1):(1'h0)]));
          reg838 = ((($unsigned($signed(forvar829)) ?
                      $signed($unsigned((8'h9c))) : reg811) ?
                  $signed((-$unsigned(reg808))) : (wire819[(3'h6):(3'h6)] * ($unsigned(reg807) ?
                      reg837[(4'hb):(3'h5)] : $signed((8'h9c))))) ?
              (+(((+forvar834) && (~wire799)) ?
                  ((reg804 ?
                      reg801 : (7'h44)) << reg804[(2'h2):(1'h1)]) : (reg806[(3'h7):(1'h0)] ?
                      $unsigned(reg807) : reg832))) : $signed(reg811[(1'h0):(1'h0)]));
          reg839 <= ((!$unsigned({(reg804 | forvar834), $signed((8'hbf))})) ?
              (reg815[(4'hd):(4'h8)] ?
                  ((reg804 ? (-reg817) : $unsigned(reg828)) ?
                      (reg832[(2'h2):(1'h1)] ?
                          (reg820 ?
                              reg838 : reg823) : $signed(reg830)) : reg800[(4'h8):(3'h4)]) : reg806) : $signed({$unsigned(reg832[(3'h4):(1'h0)])}));
        end
      reg840 <= ($unsigned(reg838) ?
          ((~&forvar834) ^ reg802) : (((reg801[(3'h7):(3'h7)] ^ ((8'haf) ?
                  reg817 : (8'ha4))) >= (&((8'hb1) != reg801))) ?
              $unsigned(forvar803) : $signed(reg833)));
      for (forvar841 = (1'h0); (forvar841 < (1'h1)); forvar841 = (forvar841 + (1'h1)))
        begin
          reg842 <= $unsigned(wire798);
          reg843 <= (~^reg818);
        end
      reg844 = reg815[(3'h7):(2'h3)];
    end
  assign wire845 = ($unsigned(reg818) ?
                       reg836[(3'h4):(2'h3)] : forvar812[(4'h8):(3'h6)]);
  module846 modinst1378 (.wire847(wire845), .y(wire1377), .wire849(reg830), .wire848(forvar834), .clk(clk), .wire850(reg804));
  always
    @(posedge clk) begin
      reg1379 <= ((^{$signed($unsigned(reg800)), {$unsigned(wire797)}}) ?
          reg816 : $signed($signed((~^$unsigned(forvar803)))));
      for (forvar1380 = (1'h0); (forvar1380 < (2'h3)); forvar1380 = (forvar1380 + (1'h1)))
        begin
          for (forvar1381 = (1'h0); (forvar1381 < (1'h0)); forvar1381 = (forvar1381 + (1'h1)))
            begin
              reg1382 = reg805;
              reg1383 <= (((reg843 ^ reg839[(3'h5):(2'h3)]) ?
                  ($signed((reg817 >> reg832)) | (^(8'hb2))) : {reg823,
                      (^{(8'ha1)})}) < ((|reg806) ?
                  {($signed((8'haf)) > (+reg818)),
                      {$unsigned(reg837)}} : ($unsigned($signed(reg823)) <<< (~^(8'ha7)))));
            end
          reg1384 <= (-$unsigned($unsigned(((^forvar821) ^~ $signed(reg800)))));
          if ((^~reg816))
            begin
              reg1385 = $unsigned($signed({(~^reg1379), wire799}));
              reg1386 = (8'hbf);
              reg1387 <= reg808[(4'ha):(4'ha)];
              reg1388 <= (((((~&reg844) ?
                              $signed(reg816) : reg833[(1'h1):(1'h1)]) ?
                          ($unsigned(reg839) << ((7'h41) ?
                              reg830 : (8'hbb))) : ({forvar1380} ?
                              reg809[(4'ha):(1'h0)] : (reg808 ?
                                  reg817 : wire1377))) ?
                      (-($unsigned(reg824) < $signed(wire798))) : ($signed(reg808[(1'h0):(1'h0)]) >>> $signed($unsigned(reg807)))) ?
                  {forvar841} : $signed((8'hac)));
            end
          else
            begin
              reg1385 = $unsigned($signed({((reg807 & (8'hbc)) <<< (8'hbc))}));
            end
          if (wire796[(1'h0):(1'h0)])
            begin
              reg1389 <= (({wire797, forvar1381} ?
                  $signed((~&reg844[(1'h0):(1'h0)])) : forvar829) * {(~^reg836[(4'hb):(4'h8)]),
                  reg833[(2'h2):(1'h1)]});
              reg1390 = wire819[(2'h3):(1'h1)];
              reg1391 = $signed((($unsigned($unsigned(wire819)) + ($unsigned(reg824) > $signed(reg831))) - reg1382));
              reg1392 <= $unsigned($signed((((7'h40) ?
                  wire810 : (wire797 - (8'hae))) - $signed((wire797 ?
                  reg806 : forvar834)))));
              reg1393 <= ((~^{(7'h42)}) ?
                  (7'h41) : $unsigned((($unsigned(reg800) ?
                      {wire798,
                          reg830} : $unsigned(forvar834)) <= (~^$signed(forvar803)))));
            end
          else
            begin
              reg1389 <= ((^reg802[(2'h3):(1'h0)]) ~^ reg1379);
              reg1390 <= reg824;
              reg1391 <= (8'hac);
            end
          reg1394 <= reg1393;
        end
      for (forvar1395 = (1'h0); (forvar1395 < (3'h4)); forvar1395 = (forvar1395 + (1'h1)))
        begin
          reg1396 <= (8'had);
        end
      reg1397 = $signed(($unsigned((-$unsigned(reg807))) ?
          $unsigned((-reg836[(5'h12):(2'h2)])) : {(!reg828)}));
      reg1398 <= reg800[(1'h0):(1'h0)];
    end
  assign wire1399 = {($unsigned((wire1377 - (wire845 ^~ (8'hb2)))) ?
                            $unsigned(($unsigned(forvar829) >> (~|wire810))) : $unsigned($signed({forvar803})))};
  assign wire1400 = $unsigned((^~((8'hb6) ?
                        {$unsigned(reg811),
                            (~reg1386)} : reg824[(2'h3):(1'h1)])));
  assign wire1401 = ((($signed($signed(reg804)) >> (8'ha8)) || (^~(reg831 ?
                        $signed((8'hba)) : (+reg1383)))) ^~ (({(reg1379 ?
                            reg1384 : (7'h40))} <= reg824[(2'h2):(1'h0)]) ^~ ((8'h9c) ^~ $signed($unsigned(reg831)))));
  always
    @(posedge clk) begin
      reg1402 = $unsigned($signed((reg806 ?
          {(forvar841 ? reg814 : reg1387)} : reg839[(2'h3):(2'h2)])));
      for (forvar1403 = (1'h0); (forvar1403 < (1'h0)); forvar1403 = (forvar1403 + (1'h1)))
        begin
          if (($signed($unsigned((|$unsigned(reg816)))) ?
              $signed((-reg809)) : {(!reg807[(3'h4):(1'h0)]),
                  reg817[(1'h1):(1'h1)]}))
            begin
              reg1404 <= forvar1403[(3'h6):(3'h4)];
            end
          else
            begin
              reg1404 <= forvar1395;
            end
        end
    end
  always
    @(posedge clk) begin
      reg1405 <= {(reg806[(1'h0):(1'h0)] ?
              ({$unsigned(reg1397), reg1386[(1'h0):(1'h0)]} ?
                  (~|(reg806 ?
                      reg1394 : wire797)) : (~$signed(reg827))) : forvar1380[(2'h2):(2'h2)])};
      reg1406 <= $signed((~|wire796[(2'h2):(1'h0)]));
      for (forvar1407 = (1'h0); (forvar1407 < (1'h1)); forvar1407 = (forvar1407 + (1'h1)))
        begin
          reg1408 <= reg1396[(3'h4):(2'h3)];
          reg1409 = $unsigned($unsigned(((reg1402[(2'h3):(2'h2)] ?
                  (8'ha9) : {reg805, reg1396}) ?
              {(reg1405 ? reg1382 : reg830),
                  (-wire819)} : $signed((reg831 ~^ reg1402)))));
          for (forvar1410 = (1'h0); (forvar1410 < (1'h1)); forvar1410 = (forvar1410 + (1'h1)))
            begin
              reg1411 <= (!$unsigned((~^$signed(reg826))));
            end
          reg1412 = forvar1407[(2'h3):(2'h3)];
          reg1413 <= reg838;
        end
      reg1414 <= $signed(({$signed((reg815 ?
              reg836 : reg1406))} ~^ $signed($signed(reg1384))));
    end
  assign wire1415 = $signed(forvar1407);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module35  (y, clk, wire36, wire37, wire38, wire39);
  output wire [(32'h2b2):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h13):(1'h0)] wire36;
  input wire [(5'h15):(1'h0)] wire37;
  input wire [(4'hd):(1'h0)] wire38;
  input wire [(3'h6):(1'h0)] wire39;
  reg [(3'h4):(1'h0)] reg786 = (1'h0);
  reg [(5'h14):(1'h0)] reg785 = (1'h0);
  reg [(4'ha):(1'h0)] reg784 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire40;
  reg signed [(5'h15):(1'h0)] reg41 = (1'h0);
  reg [(5'h12):(1'h0)] reg42 = (1'h0);
  wire [(4'hd):(1'h0)] wire162;
  wire signed [(5'h13):(1'h0)] wire164;
  wire [(5'h11):(1'h0)] wire165;
  reg signed [(3'h5):(1'h0)] forvar166 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg167 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg168 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg169 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg170 = (1'h0);
  reg [(5'h13):(1'h0)] reg171 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire172;
  wire [(4'hd):(1'h0)] wire489;
  reg [(5'h11):(1'h0)] reg491 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg492 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg493 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg494 = (1'h0);
  reg [(5'h10):(1'h0)] reg495 = (1'h0);
  reg [(3'h6):(1'h0)] forvar496 = (1'h0);
  reg [(5'h13):(1'h0)] reg497 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg498 = (1'h0);
  reg [(3'h4):(1'h0)] reg499 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg500 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg501 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg502 = (1'h0);
  reg [(5'h11):(1'h0)] reg503 = (1'h0);
  reg [(5'h13):(1'h0)] reg504 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg505 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg506 = (1'h0);
  reg [(5'h15):(1'h0)] reg507 = (1'h0);
  reg [(4'hb):(1'h0)] reg508 = (1'h0);
  wire [(3'h7):(1'h0)] wire509;
  wire signed [(5'h11):(1'h0)] wire510;
  reg signed [(4'he):(1'h0)] reg511 = (1'h0);
  reg [(5'h12):(1'h0)] reg512 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg513 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg514 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg515 = (1'h0);
  reg [(5'h13):(1'h0)] forvar516 = (1'h0);
  reg [(4'hb):(1'h0)] reg517 = (1'h0);
  reg [(3'h4):(1'h0)] reg518 = (1'h0);
  wire signed [(4'he):(1'h0)] wire519;
  wire signed [(4'he):(1'h0)] wire520;
  reg signed [(5'h13):(1'h0)] reg521 = (1'h0);
  reg [(4'hf):(1'h0)] reg522 = (1'h0);
  wire [(4'h8):(1'h0)] wire523;
  wire signed [(5'h12):(1'h0)] wire524;
  wire signed [(5'h13):(1'h0)] wire782;
  assign y = {reg786,
                 reg785,
                 reg784,
                 wire40,
                 reg41,
                 reg42,
                 wire162,
                 wire164,
                 wire165,
                 forvar166,
                 reg167,
                 reg168,
                 reg169,
                 reg170,
                 reg171,
                 wire172,
                 wire489,
                 reg491,
                 reg492,
                 reg493,
                 reg494,
                 reg495,
                 forvar496,
                 reg497,
                 reg498,
                 reg499,
                 reg500,
                 reg501,
                 reg502,
                 reg503,
                 reg504,
                 reg505,
                 reg506,
                 reg507,
                 reg508,
                 wire509,
                 wire510,
                 reg511,
                 reg512,
                 reg513,
                 reg514,
                 reg515,
                 forvar516,
                 reg517,
                 reg518,
                 wire519,
                 wire520,
                 reg521,
                 reg522,
                 wire523,
                 wire524,
                 wire782,
                 (1'h0)};
  assign wire40 = (~|{$signed($signed(((7'h44) ? wire37 : (8'hb3))))});
  always
    @(posedge clk) begin
      reg41 = ((8'haf) ~^ wire38[(3'h7):(3'h6)]);
      reg42 <= $signed(($signed($unsigned((wire39 ? (8'hb2) : reg41))) ?
          ($signed($signed(wire36)) ?
              {(wire37 ^ wire40)} : ({wire39} << reg41)) : $unsigned((^(~^wire38)))));
    end
  module43 modinst163 (.y(wire162), .wire47(wire36), .clk(clk), .wire45(wire37), .wire44(wire40), .wire46(wire38));
  assign wire164 = (+{({$signed(wire36)} * wire38)});
  assign wire165 = (8'hb7);
  always
    @(posedge clk) begin
      for (forvar166 = (1'h0); (forvar166 < (3'h4)); forvar166 = (forvar166 + (1'h1)))
        begin
          reg167 = reg41;
          reg168 <= $unsigned(wire164[(4'h8):(1'h0)]);
          reg169 <= (+(!$signed($signed((wire39 ~^ reg42)))));
          reg170 <= $signed($unsigned(({(wire164 ? wire164 : wire40),
              (wire38 || forvar166)} || $unsigned(reg41))));
          reg171 <= $unsigned(wire36);
        end
    end
  assign wire172 = (^~$unsigned((^~wire165[(3'h5):(3'h5)])));
  module173 modinst490 (.y(wire489), .wire177(reg169), .wire175(reg42), .wire174(reg41), .clk(clk), .wire176(wire36));
  always
    @(posedge clk) begin
      reg491 <= ($signed($unsigned(($unsigned(reg169) ?
          (|reg169) : $signed(wire164)))) - wire165[(4'h8):(3'h6)]);
      reg492 = ((wire162[(4'hb):(2'h3)] | wire40[(3'h5):(1'h0)]) ?
          (~(7'h44)) : $signed({(!(~wire39)), reg168[(1'h1):(1'h1)]}));
      reg493 <= $signed(($unsigned(reg491) ?
          reg41 : {(~$unsigned(forvar166)), (~$unsigned(wire37))}));
    end
  always
    @(posedge clk) begin
      reg494 = wire37[(5'h12):(5'h10)];
      if ({$signed(wire489[(1'h1):(1'h1)]), {wire165}})
        begin
          reg495 <= ($unsigned($unsigned(((wire489 & forvar166) < ((8'hb7) > reg170)))) == (^(~|(reg170 ?
              (reg168 >> reg41) : reg169))));
          for (forvar496 = (1'h0); (forvar496 < (2'h3)); forvar496 = (forvar496 + (1'h1)))
            begin
              reg497 <= reg168[(1'h1):(1'h1)];
              reg498 <= $signed({$signed($signed((wire164 ?
                      wire38 : (8'hb6))))});
              reg499 = $signed((~&(((|reg169) & (~^reg491)) ?
                  wire37[(5'h10):(3'h6)] : $unsigned(reg41))));
              reg500 <= ($unsigned($unsigned($unsigned(reg492[(4'h9):(2'h2)]))) && reg494[(2'h3):(1'h1)]);
              reg501 <= wire36;
            end
          reg502 = $unsigned(({reg42[(4'hc):(4'h8)]} ?
              (forvar166 > $unsigned(wire36)) : wire38));
          reg503 = forvar166[(3'h4):(1'h0)];
        end
      else
        begin
          reg495 <= wire172;
        end
      reg504 = (&reg491[(3'h7):(1'h1)]);
      reg505 <= reg495[(4'hf):(1'h0)];
      reg506 <= reg167;
    end
  always
    @(posedge clk) begin
      reg507 <= $signed(reg502[(3'h5):(2'h3)]);
      reg508 <= (^~(((~(wire40 ?
          wire165 : reg505)) < $signed((~wire489))) ^ ({(reg507 <<< reg167)} >>> $signed((reg499 ?
          wire165 : reg501)))));
    end
  assign wire509 = reg508[(3'h7):(2'h3)];
  assign wire510 = $signed(((reg167[(4'he):(2'h2)] ?
                           (((8'hb0) >>> reg499) ?
                               wire164 : (~&reg42)) : $signed($unsigned(reg170))) ?
                       $unsigned((wire162 > (wire489 == wire40))) : $signed((reg504[(3'h6):(1'h0)] > wire37[(1'h1):(1'h0)]))));
  always
    @(posedge clk) begin
      reg511 <= wire164;
      reg512 <= (reg492 ?
          {wire37[(4'hc):(1'h1)], reg41[(4'hf):(2'h3)]} : reg506);
      reg513 <= (!($unsigned(((^reg167) ^~ $unsigned(reg511))) | (8'hb4)));
    end
  always
    @(posedge clk) begin
      reg514 <= $signed((($unsigned((reg167 ?
              reg41 : wire40)) << ((!reg493) >>> reg494)) ?
          ($unsigned({reg508}) ? (~^(-(8'ha2))) : wire489) : reg494));
      reg515 <= reg501;
      for (forvar516 = (1'h0); (forvar516 < (1'h1)); forvar516 = (forvar516 + (1'h1)))
        begin
          reg517 <= {({(+$signed(wire165)),
                      ($unsigned(reg503) ?
                          (~reg495) : ((8'ha5) ? (8'ha5) : reg513))} ?
                  (reg41[(4'h8):(1'h0)] ?
                      reg506 : (~^$signed(wire36))) : ($unsigned(((8'hbc) || reg511)) ?
                      forvar166[(2'h3):(2'h3)] : ((-wire39) ~^ $signed(reg498)))),
              reg504[(4'hb):(3'h4)]};
          reg518 <= $unsigned($unsigned((&$signed((~reg513)))));
        end
    end
  assign wire519 = ((~&reg168[(1'h0):(1'h0)]) | $unsigned($signed((8'hbf))));
  assign wire520 = ((~$unsigned((8'ha2))) && {($unsigned(reg501[(4'hf):(4'hd)]) ?
                           ((reg502 != reg168) ~^ (~&wire489)) : (!{reg492,
                               reg500})),
                       {{{(8'hba), (8'ha1)}, (wire509 >> reg171)},
                           ((-reg517) || (reg508 ^~ wire37))}});
  always
    @(posedge clk) begin
      reg521 <= reg501[(4'hb):(2'h2)];
      reg522 <= reg501;
    end
  assign wire523 = (-$unsigned(reg513[(2'h3):(1'h1)]));
  assign wire524 = ((reg503 ?
                           $signed($unsigned((reg507 ?
                               reg168 : reg168))) : $unsigned(reg500)) ?
                       (^~reg491) : {((wire489 ?
                               reg522 : reg494[(2'h2):(2'h2)]) >= $signed(((8'hbb) < wire520)))});
  module525 modinst783 (.wire528(reg503), .wire527(wire165), .y(wire782), .wire530(wire489), .clk(clk), .wire529(reg494), .wire526(reg507));
  always
    @(posedge clk) begin
      reg784 <= ((-reg522) ?
          ((-$unsigned(reg514)) + (!((^~(8'hba)) ?
              {(8'hb4)} : wire520))) : $signed($signed(reg167[(2'h3):(1'h0)])));
      reg785 = {reg505[(2'h2):(2'h2)]};
      reg786 <= (wire782[(5'h13):(5'h10)] > $signed($unsigned((((8'ha3) ?
              wire165 : reg785) ?
          $signed((7'h40)) : wire782))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module525
#(parameter param781 = (8'hbb))
(y, clk, wire530, wire529, wire528, wire527, wire526);
  output wire [(32'h348):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire530;
  input wire [(4'h8):(1'h0)] wire529;
  input wire [(5'h11):(1'h0)] wire528;
  input wire signed [(5'h10):(1'h0)] wire527;
  input wire [(5'h15):(1'h0)] wire526;
  wire signed [(4'h8):(1'h0)] wire780;
  reg [(4'h9):(1'h0)] reg779 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg765 = (1'h0);
  reg [(4'hd):(1'h0)] reg778 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg777 = (1'h0);
  reg [(3'h7):(1'h0)] reg776 = (1'h0);
  reg [(4'hc):(1'h0)] reg775 = (1'h0);
  reg [(4'hf):(1'h0)] reg774 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg773 = (1'h0);
  reg [(5'h11):(1'h0)] forvar772 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg771 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg770 = (1'h0);
  reg [(5'h15):(1'h0)] reg769 = (1'h0);
  reg [(5'h13):(1'h0)] reg768 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg767 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg766 = (1'h0);
  reg [(4'hc):(1'h0)] forvar765 = (1'h0);
  reg [(4'hd):(1'h0)] reg764 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg763 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg762 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar761 = (1'h0);
  reg [(5'h13):(1'h0)] forvar760 = (1'h0);
  reg [(4'ha):(1'h0)] reg759 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg758 = (1'h0);
  reg [(4'hb):(1'h0)] reg757 = (1'h0);
  reg [(4'hb):(1'h0)] reg756 = (1'h0);
  wire [(5'h10):(1'h0)] wire649;
  reg [(5'h15):(1'h0)] reg532 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg531 = (1'h0);
  reg [(4'he):(1'h0)] reg651 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg652 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg653 = (1'h0);
  reg [(3'h7):(1'h0)] reg654 = (1'h0);
  reg [(3'h4):(1'h0)] forvar655 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg656 = (1'h0);
  reg [(3'h6):(1'h0)] forvar657 = (1'h0);
  reg [(2'h3):(1'h0)] reg658 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg659 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg660 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg661 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg662 = (1'h0);
  reg [(5'h14):(1'h0)] reg663 = (1'h0);
  reg [(3'h4):(1'h0)] reg664 = (1'h0);
  reg [(4'h8):(1'h0)] reg665 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg666 = (1'h0);
  reg [(4'hd):(1'h0)] reg667 = (1'h0);
  reg [(3'h7):(1'h0)] reg668 = (1'h0);
  reg signed [(4'he):(1'h0)] reg669 = (1'h0);
  reg [(4'hc):(1'h0)] reg670 = (1'h0);
  reg [(4'he):(1'h0)] forvar671 = (1'h0);
  reg [(5'h12):(1'h0)] reg672 = (1'h0);
  reg [(4'h9):(1'h0)] reg673 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg674 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg675 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg676 = (1'h0);
  reg [(5'h12):(1'h0)] reg677 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg678 = (1'h0);
  reg [(2'h3):(1'h0)] reg679 = (1'h0);
  reg [(4'hf):(1'h0)] reg680 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg681 = (1'h0);
  reg [(3'h7):(1'h0)] reg682 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg683 = (1'h0);
  reg [(3'h5):(1'h0)] reg684 = (1'h0);
  reg [(3'h5):(1'h0)] reg685 = (1'h0);
  reg [(3'h5):(1'h0)] reg686 = (1'h0);
  reg [(4'h9):(1'h0)] reg687 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire754;
  assign y = {wire780,
                 reg779,
                 reg765,
                 reg778,
                 reg777,
                 reg776,
                 reg775,
                 reg774,
                 reg773,
                 forvar772,
                 reg771,
                 reg770,
                 reg769,
                 reg768,
                 reg767,
                 reg766,
                 forvar765,
                 reg764,
                 reg763,
                 reg762,
                 forvar761,
                 forvar760,
                 reg759,
                 reg758,
                 reg757,
                 reg756,
                 wire649,
                 reg532,
                 reg531,
                 reg651,
                 reg652,
                 reg653,
                 reg654,
                 forvar655,
                 reg656,
                 forvar657,
                 reg658,
                 reg659,
                 reg660,
                 reg661,
                 reg662,
                 reg663,
                 reg664,
                 reg665,
                 reg666,
                 reg667,
                 reg668,
                 reg669,
                 reg670,
                 forvar671,
                 reg672,
                 reg673,
                 reg674,
                 reg675,
                 reg676,
                 reg677,
                 reg678,
                 reg679,
                 reg680,
                 reg681,
                 reg682,
                 reg683,
                 reg684,
                 reg685,
                 reg686,
                 reg687,
                 wire754,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg531 = $signed(wire529[(4'h8):(3'h7)]);
      reg532 = $unsigned((^$signed(wire528)));
    end
  module533 modinst650 (.wire536(wire526), .clk(clk), .wire538(wire527), .wire534(wire528), .wire537(wire530), .wire535(reg531), .y(wire649));
  always
    @(posedge clk) begin
      reg651 = (wire526[(5'h13):(4'h8)] <<< wire527);
    end
  always
    @(posedge clk) begin
      reg652 <= {$signed(wire527), wire526};
      reg653 = wire530[(4'h9):(3'h7)];
      reg654 <= ($signed(wire530[(4'h9):(1'h0)]) <= (wire649[(5'h10):(3'h4)] ?
          $unsigned(reg652) : (((~wire527) ?
                  (~reg531) : wire649[(4'hb):(4'h9)]) ?
              $unsigned((reg652 && wire526)) : {wire649, reg531})));
      for (forvar655 = (1'h0); (forvar655 < (2'h3)); forvar655 = (forvar655 + (1'h1)))
        begin
          reg656 = reg654;
          for (forvar657 = (1'h0); (forvar657 < (1'h0)); forvar657 = (forvar657 + (1'h1)))
            begin
              reg658 = (~|(~wire527[(1'h1):(1'h1)]));
              reg659 <= reg658;
              reg660 <= (8'hb3);
            end
          reg661 = $unsigned((reg653 ?
              reg659 : $unsigned(((forvar657 >>> wire649) < (~&wire528)))));
          reg662 <= (&(+wire527[(2'h2):(1'h0)]));
          reg663 <= $signed(($signed(wire527[(4'hc):(1'h1)]) ?
              $signed(($signed(wire526) | (reg662 > reg662))) : (8'hb1)));
        end
    end
  always
    @(posedge clk) begin
      reg664 <= $signed((~^$unsigned(reg659[(1'h1):(1'h1)])));
      reg665 <= $unsigned($signed($signed(reg664[(2'h2):(1'h1)])));
    end
  always
    @(posedge clk) begin
      reg666 <= reg663;
      reg667 = (|$signed((8'ha1)));
      reg668 <= (reg660[(4'h9):(3'h5)] ?
          $signed((!reg651)) : reg658[(2'h3):(2'h3)]);
    end
  always
    @(posedge clk) begin
      reg669 <= ($signed($signed($unsigned((7'h44)))) >>> $signed(reg660[(4'h8):(3'h4)]));
      reg670 <= reg652;
      for (forvar671 = (1'h0); (forvar671 < (3'h4)); forvar671 = (forvar671 + (1'h1)))
        begin
          reg672 <= {((reg667[(3'h7):(3'h6)] <= $unsigned(reg654[(2'h3):(1'h1)])) || forvar671[(4'ha):(4'h8)])};
          reg673 <= $signed(((~^reg668[(1'h1):(1'h1)]) > $signed(reg661[(2'h3):(1'h0)])));
          reg674 <= $signed((wire649 ?
              $signed($signed((reg665 ?
                  reg653 : reg651))) : (+(+reg660[(5'h13):(4'he)]))));
          reg675 = reg665;
          reg676 <= $unsigned((reg660 ? reg656[(2'h3):(1'h0)] : reg670));
        end
      reg677 <= (reg674[(3'h5):(2'h3)] ?
          ({(reg656[(2'h3):(2'h2)] & reg667)} ?
              (reg652 & (forvar657[(3'h4):(1'h1)] ?
                  (reg661 == reg664) : (reg662 ?
                      reg666 : reg662))) : (((forvar657 ^ forvar655) && wire649[(4'hd):(1'h1)]) ?
                  $signed((reg663 ~^ reg674)) : ((~&forvar657) >>> ((8'hb9) > reg672)))) : ($signed(forvar655[(1'h1):(1'h0)]) ?
              reg663[(4'hd):(3'h6)] : reg653[(3'h4):(1'h0)]));
    end
  always
    @(posedge clk) begin
      reg678 = (!((!forvar671[(4'h8):(3'h6)]) ?
          (|$unsigned($signed(wire530))) : $signed(reg665)));
      reg679 = (wire649[(3'h6):(3'h5)] ?
          $signed((reg678 ?
              (&(reg670 && reg661)) : ($unsigned(wire529) || (~&wire529)))) : reg672);
      reg680 <= $signed((-($signed(reg656) ? {$signed(reg677)} : wire529)));
      reg681 <= {reg672[(4'hf):(4'hb)]};
      reg682 <= $signed(reg675);
    end
  always
    @(posedge clk) begin
      reg683 <= ($unsigned((((-reg660) ?
                  (reg532 ? wire527 : (8'h9f)) : reg665) ?
              {$signed(wire528), $signed(reg669)} : reg661)) ?
          (((~(forvar655 || reg651)) && $signed((~^wire528))) < wire526[(4'ha):(2'h3)]) : (~|reg665[(3'h5):(1'h0)]));
      reg684 <= ((reg669[(1'h1):(1'h0)] ?
          (reg656 ?
              (~|$signed(reg669)) : (8'hb6)) : $unsigned(((reg681 & reg670) ~^ {reg532,
              (8'ha0)}))) & $signed((~wire530[(3'h7):(2'h2)])));
      reg685 <= {reg651[(3'h6):(1'h0)]};
      reg686 <= $unsigned(($signed(forvar671) ?
          $unsigned(((8'hb9) ? ((8'hab) + (7'h43)) : reg663)) : reg681));
      reg687 = ((reg680 >>> {{$unsigned(forvar671)}}) ?
          $unsigned($unsigned(reg669)) : $signed((^{reg670[(3'h5):(2'h2)],
              $signed(reg662)})));
    end
  module688 modinst755 (wire754, clk, reg670, reg674, reg652, reg683, reg661);
  always
    @(posedge clk) begin
      reg756 <= forvar671;
      reg757 <= ((~^(~&reg661[(4'hc):(4'h9)])) != $unsigned((-(forvar671[(4'h9):(3'h6)] <<< (reg681 <= reg651)))));
      reg758 <= reg656[(2'h3):(2'h3)];
    end
  always
    @(posedge clk) begin
      reg759 <= $unsigned((+(!(8'had))));
    end
  always
    @(posedge clk) begin
      for (forvar760 = (1'h0); (forvar760 < (1'h1)); forvar760 = (forvar760 + (1'h1)))
        begin
          for (forvar761 = (1'h0); (forvar761 < (1'h1)); forvar761 = (forvar761 + (1'h1)))
            begin
              reg762 <= $signed(((+reg685) <= {$signed((reg685 <= reg676))}));
            end
          reg763 <= (reg687 ^~ $unsigned((reg687 & (8'ha7))));
        end
      reg764 = (~(reg662[(3'h7):(1'h1)] ?
          (|reg662) : ((~&$signed(reg665)) ? reg759[(3'h6):(3'h5)] : reg757)));
      if ((^(reg686[(3'h5):(1'h1)] <= (^reg680))))
        begin
          for (forvar765 = (1'h0); (forvar765 < (1'h0)); forvar765 = (forvar765 + (1'h1)))
            begin
              reg766 = ({{wire529,
                      $unsigned((~|reg532))}} < reg680[(2'h3):(2'h3)]);
              reg767 <= (((+(~|wire527[(2'h2):(1'h1)])) ?
                      ({$signed(wire754),
                          (|(8'hb5))} >>> reg682[(1'h1):(1'h0)]) : (8'hb5)) ?
                  (-wire526) : reg532[(4'hc):(4'h8)]);
              reg768 <= (~|(reg674[(4'ha):(3'h7)] ?
                  (^~wire649[(4'he):(3'h5)]) : $signed(($signed(wire649) ~^ (reg762 ?
                      reg673 : reg654)))));
              reg769 <= ($unsigned((($signed(wire649) ?
                          (reg679 <<< reg685) : reg759[(4'h9):(3'h6)]) ?
                      $unsigned((reg665 ? (8'hb2) : reg678)) : {$signed(reg756),
                          {reg667}})) ?
                  reg670 : reg764);
              reg770 = {reg673, {$unsigned(reg676), wire754}};
            end
          reg771 = $signed({{($signed(reg678) ?
                      (wire529 ? forvar655 : wire529) : (reg674 < forvar671)),
                  (&$unsigned(wire527))},
              reg656});
          for (forvar772 = (1'h0); (forvar772 < (1'h1)); forvar772 = (forvar772 + (1'h1)))
            begin
              reg773 <= ($signed({reg674}) >>> (&$unsigned(((reg769 ?
                  reg651 : reg675) >>> $unsigned(reg766)))));
              reg774 = (forvar655[(2'h3):(2'h2)] ?
                  ((reg654 || reg764) ?
                      $signed($signed((reg770 ? reg653 : reg680))) : (-(reg666 ?
                          reg668 : {reg659}))) : ({forvar761} ?
                      reg769 : $unsigned(forvar761[(4'h8):(2'h2)])));
              reg775 <= {(~|(+$signed((wire526 ? reg679 : wire529)))), reg674};
              reg776 = $signed((8'hb3));
              reg777 = $signed({$unsigned(((reg653 ? forvar655 : (8'hba)) ?
                      reg680 : (wire754 < wire754))),
                  $unsigned((^(reg686 ? reg663 : reg766)))});
            end
          reg778 <= $unsigned(reg674);
        end
      else
        begin
          reg765 <= ($signed(reg767[(2'h2):(1'h0)]) < ($unsigned(((+(8'hb2)) <= (reg756 ?
              reg776 : (8'h9c)))) ^~ (~&(~^(reg653 ? reg654 : (8'hac))))));
          reg766 = reg666;
          reg767 <= (^~{(((reg764 ?
                  reg775 : (8'ha9)) + reg669[(1'h0):(1'h0)]) || (|(reg776 ?
                  reg672 : reg684))),
              (~&$unsigned(reg777))});
        end
    end
  always
    @(posedge clk) begin
      reg779 <= (((($unsigned(reg680) ?
                      (reg663 ? reg654 : reg670) : $signed(forvar655)) ?
                  forvar760[(1'h1):(1'h1)] : ($unsigned(reg663) ?
                      $unsigned(reg652) : reg667)) ?
              reg771[(3'h7):(2'h2)] : $unsigned({$signed(reg659)})) ?
          (&$signed(reg682)) : $unsigned((7'h44)));
    end
  assign wire780 = reg663[(4'hc):(2'h2)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module173
#( parameter param488 = (~&((({(8'h9f)} ? ((8'hbf) ? (8'hae) : (8'hbb)) : (~(8'hab))) ? (((8'h9f) ? (8'haf) : (7'h40)) | (^(8'hbd))) : ((8'haa) ? {(8'hac), (8'hb9)} : {(8'hbe)})) ? {(((8'hab) ? (8'hb3) : (8'h9d)) ? ((8'hbf) << (8'had)) : ((8'ha9) >>> (7'h42)))} : {{((8'ha5) == (8'hbf)), ((8'hb4) <<< (8'ha6))}, {(-(8'ha6))}})) )
(y, clk, wire177, wire176, wire175, wire174);
  output wire [(32'h2b3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h12):(1'h0)] wire177;
  input wire [(5'h13):(1'h0)] wire176;
  input wire signed [(3'h5):(1'h0)] wire175;
  input wire signed [(4'ha):(1'h0)] wire174;
  reg [(3'h5):(1'h0)] reg487 = (1'h0);
  reg [(5'h12):(1'h0)] reg486 = (1'h0);
  reg [(2'h2):(1'h0)] reg485 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg484 = (1'h0);
  reg [(4'h9):(1'h0)] reg483 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg482 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg481 = (1'h0);
  reg [(3'h5):(1'h0)] reg480 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar479 = (1'h0);
  reg [(3'h7):(1'h0)] reg478 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar477 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg476 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg475 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg474 = (1'h0);
  reg [(5'h14):(1'h0)] forvar473 = (1'h0);
  reg [(3'h4):(1'h0)] reg472 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar471 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire470;
  reg signed [(5'h11):(1'h0)] reg469 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg468 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg467 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg466 = (1'h0);
  reg [(5'h10):(1'h0)] reg465 = (1'h0);
  reg signed [(4'he):(1'h0)] reg464 = (1'h0);
  reg [(5'h11):(1'h0)] reg463 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire462;
  wire [(4'hf):(1'h0)] wire460;
  reg [(2'h3):(1'h0)] reg212 = (1'h0);
  reg [(5'h13):(1'h0)] reg211 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar210 = (1'h0);
  reg [(5'h10):(1'h0)] reg209 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg208 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar207 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg206 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg205 = (1'h0);
  reg [(4'hb):(1'h0)] reg204 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire203;
  reg [(4'h9):(1'h0)] reg202 = (1'h0);
  reg [(4'hc):(1'h0)] reg201 = (1'h0);
  reg [(4'he):(1'h0)] reg200 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg199 = (1'h0);
  reg [(4'h9):(1'h0)] reg191 = (1'h0);
  reg [(3'h4):(1'h0)] reg198 = (1'h0);
  reg [(4'h8):(1'h0)] reg197 = (1'h0);
  reg [(3'h7):(1'h0)] forvar196 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg195 = (1'h0);
  reg [(4'h9):(1'h0)] reg194 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg193 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg192 = (1'h0);
  reg [(4'hd):(1'h0)] forvar191 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg190 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire189;
  wire signed [(4'h9):(1'h0)] wire188;
  wire signed [(5'h12):(1'h0)] wire187;
  reg [(4'he):(1'h0)] reg186 = (1'h0);
  reg [(3'h4):(1'h0)] reg185 = (1'h0);
  reg [(5'h14):(1'h0)] reg184 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar183 = (1'h0);
  reg [(4'h9):(1'h0)] reg182 = (1'h0);
  reg [(5'h10):(1'h0)] reg181 = (1'h0);
  reg signed [(4'he):(1'h0)] reg180 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg179 = (1'h0);
  wire [(3'h4):(1'h0)] wire178;
  assign y = {reg487,
                 reg486,
                 reg485,
                 reg484,
                 reg483,
                 reg482,
                 reg481,
                 reg480,
                 forvar479,
                 reg478,
                 forvar477,
                 reg476,
                 reg475,
                 reg474,
                 forvar473,
                 reg472,
                 forvar471,
                 wire470,
                 reg469,
                 reg468,
                 reg467,
                 reg466,
                 reg465,
                 reg464,
                 reg463,
                 wire462,
                 wire460,
                 reg212,
                 reg211,
                 forvar210,
                 reg209,
                 reg208,
                 forvar207,
                 reg206,
                 reg205,
                 reg204,
                 wire203,
                 reg202,
                 reg201,
                 reg200,
                 reg199,
                 reg191,
                 reg198,
                 reg197,
                 forvar196,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 forvar191,
                 reg190,
                 wire189,
                 wire188,
                 wire187,
                 reg186,
                 reg185,
                 reg184,
                 forvar183,
                 reg182,
                 reg181,
                 reg180,
                 reg179,
                 wire178,
                 (1'h0)};
  assign wire178 = $unsigned(((~^{{wire174}}) || wire174[(3'h5):(1'h1)]));
  always
    @(posedge clk) begin
      reg179 = ((~^{wire177[(4'h8):(3'h6)],
          wire175[(3'h4):(3'h4)]}) | $unsigned(wire178));
      reg180 = $signed({(~|(~$signed(wire177))),
          $unsigned($unsigned($unsigned(wire176)))});
      reg181 <= ((wire178[(1'h1):(1'h0)] ?
          (reg180 ?
              $signed($signed(wire175)) : ($signed(reg180) ?
                  wire176 : reg180)) : reg180) - {((~|{reg180}) < reg180)});
    end
  always
    @(posedge clk) begin
      reg182 = {(((|$unsigned((8'haf))) ? wire175 : $unsigned(wire177)) ?
              (~&wire175[(3'h5):(3'h4)]) : ((-(&reg181)) && ({(7'h42), reg181} ?
                  $unsigned(reg181) : $unsigned(wire177))))};
      for (forvar183 = (1'h0); (forvar183 < (2'h3)); forvar183 = (forvar183 + (1'h1)))
        begin
          reg184 = $signed($signed((((~|reg182) <<< reg180[(3'h5):(2'h2)]) ?
              wire177[(4'h9):(3'h5)] : {(wire176 ? wire176 : wire177)})));
          reg185 <= $signed((wire174 ?
              wire174[(4'ha):(3'h7)] : wire178[(2'h3):(2'h2)]));
        end
      reg186 <= (~&(wire176 ?
          ((|$unsigned(reg182)) ?
              ((wire174 ^~ reg185) || $signed(reg182)) : (~|$signed(wire177))) : (|($signed(reg184) ?
              reg180[(4'ha):(1'h1)] : wire178))));
    end
  assign wire187 = (wire178[(1'h0):(1'h0)] ~^ ($unsigned($unsigned((wire178 <= reg184))) << (~^$signed(forvar183[(3'h6):(2'h2)]))));
  assign wire188 = $unsigned((reg186[(1'h1):(1'h1)] ?
                       $unsigned(wire174[(2'h2):(2'h2)]) : reg185[(3'h4):(3'h4)]));
  assign wire189 = (8'ha5);
  always
    @(posedge clk) begin
      if ($signed(reg181[(2'h2):(1'h0)]))
        begin
          reg190 = $signed(wire176[(1'h1):(1'h0)]);
          for (forvar191 = (1'h0); (forvar191 < (3'h4)); forvar191 = (forvar191 + (1'h1)))
            begin
              reg192 <= (((~|(~^(reg180 >= reg181))) >>> $unsigned(reg182)) >= reg186[(4'he):(2'h3)]);
              reg193 <= ({reg185} ?
                  wire187[(3'h7):(3'h6)] : ((wire177 ?
                          wire178[(2'h2):(2'h2)] : ((wire177 ?
                                  forvar191 : reg185) ?
                              $signed(reg190) : reg190)) ?
                      (wire187 ?
                          (+wire174[(3'h7):(1'h1)]) : ((reg186 || reg180) ?
                              (!reg192) : {(8'hbf)})) : $signed(((reg184 >> wire188) ?
                          (wire187 ?
                              forvar191 : reg184) : (reg179 < wire187)))));
              reg194 <= ($unsigned($signed(reg182[(1'h1):(1'h1)])) ?
                  forvar191 : ((^$signed(wire188[(4'h8):(3'h6)])) | ((~(~&reg179)) >= (~wire175[(2'h2):(2'h2)]))));
            end
          reg195 <= $signed({$signed($unsigned(reg182[(4'h8):(4'h8)])),
              forvar183[(3'h4):(2'h2)]});
          for (forvar196 = (1'h0); (forvar196 < (3'h4)); forvar196 = (forvar196 + (1'h1)))
            begin
              reg197 <= (((~(~^wire189)) + (!$unsigned((|reg194)))) != (reg185[(1'h0):(1'h0)] ?
                  reg184 : ($unsigned((forvar183 | reg192)) ?
                      {(forvar196 ? reg179 : reg179),
                          (reg180 ? reg181 : wire188)} : $signed((|wire189)))));
            end
          reg198 <= (wire189 >= $unsigned((&$signed((8'ha3)))));
        end
      else
        begin
          reg190 <= reg197[(2'h2):(1'h0)];
          reg191 <= {(+forvar191)};
          reg192 = $signed(({reg184[(1'h0):(1'h0)],
              $unsigned((reg195 ^~ reg192))} == $unsigned($signed(wire175))));
          reg193 = $unsigned(reg179[(1'h1):(1'h1)]);
          reg194 <= reg179;
        end
      reg199 = $signed($signed($unsigned(reg195)));
      reg200 <= (^reg197[(3'h6):(3'h4)]);
      reg201 <= $signed(({{reg182, $signed(reg186)},
          ($signed(reg181) ?
              (wire187 ?
                  (7'h43) : wire188) : $unsigned(reg184))} >>> ($signed($unsigned(wire176)) > (+((8'hb9) >> reg198)))));
    end
  always
    @(posedge clk) begin
      reg202 = ((8'h9d) < {$signed(((^~(8'hab)) ? (!wire178) : (8'haf)))});
    end
  assign wire203 = wire188[(4'h9):(4'h9)];
  always
    @(posedge clk) begin
      reg204 = ($unsigned($unsigned({$signed(forvar196),
              reg186[(3'h4):(3'h4)]})) ?
          (($signed(((8'hb8) ? wire177 : (8'ha4))) * {reg199}) ?
              $unsigned(wire188) : (-(8'hb9))) : $signed($signed(($unsigned(reg191) - (+reg200)))));
    end
  always
    @(posedge clk) begin
      reg205 = ($unsigned((^(forvar196[(3'h5):(2'h2)] ?
          forvar196 : $signed((8'h9d))))) + (~&(+reg184)));
      reg206 <= (8'hb0);
      for (forvar207 = (1'h0); (forvar207 < (1'h0)); forvar207 = (forvar207 + (1'h1)))
        begin
          reg208 <= $unsigned(((({reg180} ?
                  reg204[(4'hb):(4'h9)] : {wire176, (8'ha4)}) ?
              $unsigned((forvar196 ?
                  (8'ha3) : reg191)) : (7'h41)) <<< $unsigned(wire176[(2'h3):(1'h1)])));
          reg209 <= reg198[(3'h4):(2'h3)];
          for (forvar210 = (1'h0); (forvar210 < (1'h0)); forvar210 = (forvar210 + (1'h1)))
            begin
              reg211 <= (~^forvar183[(2'h3):(2'h2)]);
            end
          reg212 = wire188;
        end
    end
  module213 modinst461 (.wire215(wire177), .wire217(wire176), .y(wire460), .clk(clk), .wire214(reg181), .wire216(forvar210));
  assign wire462 = reg199;
  always
    @(posedge clk) begin
      reg463 = ((((!(!reg180)) ?
              reg179 : $unsigned(wire178[(1'h0):(1'h0)])) << forvar207[(4'h9):(4'h9)]) ?
          (8'h9d) : reg181);
    end
  always
    @(posedge clk) begin
      reg464 <= forvar191[(4'ha):(2'h2)];
      reg465 <= {(($signed((reg212 ? reg197 : wire174)) ?
              $signed($signed(wire189)) : wire177) * reg198)};
    end
  always
    @(posedge clk) begin
      reg466 <= (|(reg181 ?
          (reg192[(1'h0):(1'h0)] ? reg464 : (8'hb9)) : $unsigned((-((8'ha0) ?
              wire462 : reg202)))));
      reg467 = reg197[(2'h2):(1'h1)];
      reg468 <= reg190;
      reg469 = reg209;
    end
  assign wire470 = {(-((|(-wire177)) ?
                           ($signed(reg466) ?
                               {reg201} : (wire460 - reg467)) : (|reg179)))};
  always
    @(posedge clk) begin
      for (forvar471 = (1'h0); (forvar471 < (1'h1)); forvar471 = (forvar471 + (1'h1)))
        begin
          reg472 = (($unsigned(wire176) ?
              reg197[(1'h1):(1'h1)] : (~&reg465)) >= (reg197 ?
              (($signed((8'hbc)) > (wire462 ?
                  wire462 : (8'hb6))) ~^ (&(^reg467))) : (reg180[(4'hb):(1'h0)] ?
                  $signed((~&reg204)) : reg179)));
          for (forvar473 = (1'h0); (forvar473 < (3'h4)); forvar473 = (forvar473 + (1'h1)))
            begin
              reg474 = reg467;
              reg475 <= ($signed((reg201 ?
                      $signed(((8'ha7) > (8'hab))) : wire175[(2'h2):(1'h0)])) ?
                  (reg199 ?
                      $unsigned($signed((reg200 != reg474))) : (($unsigned((8'ha9)) ?
                          wire188 : (~&reg463)) && $unsigned($unsigned((8'ha1))))) : $signed((((reg464 ?
                              reg212 : (7'h44)) ?
                          reg200[(4'hc):(3'h6)] : (reg466 ? (8'ha0) : reg205)) ?
                      ((|reg469) ?
                          (~reg193) : (reg472 ?
                              forvar191 : forvar207)) : (&(reg469 ?
                          wire175 : reg180)))));
            end
          reg476 <= ({(((forvar196 ? reg465 : (8'hb4)) ? reg198 : reg212) ?
                  ($signed(reg198) ?
                      (8'ha9) : wire203) : $unsigned((reg475 - reg180)))} == {reg206[(2'h2):(1'h0)],
              ((8'ha2) >= (!{forvar207}))});
          for (forvar477 = (1'h0); (forvar477 < (2'h2)); forvar477 = (forvar477 + (1'h1)))
            begin
              reg478 <= (!$unsigned($unsigned(wire175)));
            end
          for (forvar479 = (1'h0); (forvar479 < (1'h1)); forvar479 = (forvar479 + (1'h1)))
            begin
              reg480 <= (reg191 ?
                  (^~((^$unsigned((8'hbe))) ?
                      reg192[(3'h4):(2'h3)] : (&(reg202 ?
                          wire470 : reg208)))) : $signed({reg211[(4'h9):(4'h8)]}));
              reg481 <= (&((reg463 - $signed((!wire462))) ?
                  $unsigned((8'hbd)) : (((|reg465) ?
                      (forvar207 ? reg205 : reg209) : (~|reg180)) | (forvar471 ?
                      $unsigned(reg181) : reg201))));
              reg482 = {({$unsigned((^reg475))} >> (((-wire176) * (^reg478)) + forvar196)),
                  $signed(reg472)};
              reg483 <= $unsigned((~^reg195[(1'h1):(1'h0)]));
            end
        end
      reg484 <= (reg202[(2'h2):(1'h1)] ?
          ($unsigned((|(!reg205))) ?
              {(&reg464[(3'h4):(3'h4)]), reg481} : reg211) : (8'ha1));
      reg485 <= reg193;
      reg486 <= reg469;
      reg487 <= ($unsigned((((~|reg198) ? reg466[(4'he):(3'h5)] : (~|(8'hba))) ?
          (+reg185) : {((7'h40) << reg481)})) << (+(~&(reg195[(2'h3):(1'h1)] << $unsigned(reg179)))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module43
#(parameter param161 = (8'h9c))
(y, clk, wire47, wire46, wire45, wire44);
  output wire [(32'hf6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire47;
  input wire signed [(4'ha):(1'h0)] wire46;
  input wire signed [(5'h15):(1'h0)] wire45;
  input wire [(4'ha):(1'h0)] wire44;
  reg [(3'h5):(1'h0)] reg160 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg159 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar158 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire157;
  wire signed [(4'hf):(1'h0)] wire156;
  reg [(4'he):(1'h0)] reg155 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg154 = (1'h0);
  reg [(4'ha):(1'h0)] reg153 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg152 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg151 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire149;
  wire [(5'h14):(1'h0)] wire56;
  wire signed [(4'hb):(1'h0)] wire55;
  wire [(3'h7):(1'h0)] wire54;
  reg [(5'h14):(1'h0)] reg53 = (1'h0);
  reg [(4'hc):(1'h0)] reg52 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg51 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg50 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg49 = (1'h0);
  wire [(5'h13):(1'h0)] wire48;
  assign y = {reg160,
                 reg159,
                 forvar158,
                 wire157,
                 wire156,
                 reg155,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 wire149,
                 wire56,
                 wire55,
                 wire54,
                 reg53,
                 reg52,
                 reg51,
                 reg50,
                 reg49,
                 wire48,
                 (1'h0)};
  assign wire48 = $signed($unsigned($unsigned($signed((8'hba)))));
  always
    @(posedge clk) begin
      reg49 <= {$unsigned((|{wire47[(3'h7):(2'h3)]}))};
      reg50 <= (~|$unsigned((wire45 ?
          {(^~reg49), (reg49 >>> (7'h44))} : $signed({wire47}))));
      reg51 = wire46;
    end
  always
    @(posedge clk) begin
      reg52 <= (8'hae);
      reg53 <= reg51;
    end
  assign wire54 = $unsigned($unsigned($unsigned(((~|reg50) ?
                      ((8'hb9) ? (8'hb8) : wire45) : $unsigned(wire47)))));
  assign wire55 = wire44;
  assign wire56 = wire46[(3'h7):(1'h0)];
  module57 modinst150 (wire149, clk, reg53, wire45, wire56, wire44);
  always
    @(posedge clk) begin
      reg151 <= {{$signed($signed(wire44)),
              (wire55 == (wire56[(1'h1):(1'h0)] ?
                  ((8'h9f) ? reg49 : wire56) : (~&wire48)))}};
      reg152 <= $signed(($unsigned((8'hb4)) ? (8'ha5) : reg50));
      reg153 <= (!$signed($unsigned(wire45[(5'h12):(4'he)])));
      reg154 <= (reg50[(1'h0):(1'h0)] >>> $signed((~&wire48[(1'h1):(1'h1)])));
      reg155 <= wire45;
    end
  assign wire156 = reg53;
  assign wire157 = $signed($signed((~&reg151[(1'h0):(1'h0)])));
  always
    @(posedge clk) begin
      for (forvar158 = (1'h0); (forvar158 < (2'h2)); forvar158 = (forvar158 + (1'h1)))
        begin
          reg159 = $unsigned((((&(forvar158 > forvar158)) << reg49[(4'ha):(3'h7)]) ?
              $unsigned(($signed(wire56) ?
                  ((8'h9d) ?
                      wire156 : wire47) : reg153)) : reg151[(3'h7):(1'h1)]));
          reg160 <= ($unsigned($signed({(reg50 ~^ reg153),
                  reg152[(3'h7):(3'h5)]})) ?
              ($unsigned((forvar158 >> (-(8'ha1)))) ?
                  (((~&reg49) ^ $unsigned(reg151)) >= ({reg49, wire149} ?
                      (reg152 ^ wire44) : $unsigned(reg53))) : ({$signed(reg49),
                          wire48[(1'h1):(1'h1)]} ?
                      reg51 : (reg151 ?
                          $unsigned(wire45) : (^~wire46)))) : (wire156[(4'he):(4'hc)] ^ $signed($unsigned($signed(reg52)))));
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module57
#( parameter param147 = (((^(^(~(8'hba)))) ? ((((8'haf) ^~ (8'hba)) ? (8'hab) : ((8'hb7) <<< (8'hb8))) > (((7'h40) ^~ (8'h9e)) ? {(8'hbe), (7'h44)} : ((8'hba) <<< (8'ha7)))) : ((((8'haf) <<< (8'ha0)) || (~^(8'ha7))) ? (^((8'hba) ? (8'ha7) : (8'hb9))) : (+{(8'hac), (8'h9d)}))) ? {(~^(((8'hab) ? (8'h9c) : (8'hb6)) ? ((8'hb3) - (7'h41)) : ((8'hb7) > (8'hbc))))} : (^((((8'hb1) ? (8'hb9) : (8'hb5)) ? ((8'h9d) ? (8'hb9) : (7'h40)) : ((7'h40) ? (8'hb9) : (8'hab))) ? (8'hb2) : {{(8'hb9)}})))
, parameter param148 = ({{((!(8'ha1)) ~^ (~param147))}} ? ((^~((-param147) ~^ {param147, param147})) ? param147 : {(((8'hba) ? param147 : param147) + param147), (~|(^(8'h9d)))}) : {{param147, (8'hb5)}}) )
(y, clk, wire58, wire59, wire60, wire61);
  output wire [(32'hdc):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire58;
  input wire [(4'hc):(1'h0)] wire59;
  input wire [(5'h14):(1'h0)] wire60;
  input wire signed [(2'h2):(1'h0)] wire61;
  wire [(5'h11):(1'h0)] wire146;
  wire [(5'h15):(1'h0)] wire145;
  reg [(4'hc):(1'h0)] reg144 = (1'h0);
  reg [(3'h7):(1'h0)] reg143 = (1'h0);
  reg [(4'hc):(1'h0)] reg142 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg141 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg62 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg63 = (1'h0);
  reg [(5'h12):(1'h0)] reg64 = (1'h0);
  reg [(2'h2):(1'h0)] forvar65 = (1'h0);
  reg [(4'ha):(1'h0)] reg66 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar67 = (1'h0);
  reg [(5'h14):(1'h0)] reg68 = (1'h0);
  reg [(4'ha):(1'h0)] reg69 = (1'h0);
  reg [(4'ha):(1'h0)] reg70 = (1'h0);
  reg [(2'h2):(1'h0)] reg71 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg72 = (1'h0);
  wire signed [(4'he):(1'h0)] wire139;
  assign y = {wire146,
                 wire145,
                 reg144,
                 reg143,
                 reg142,
                 reg141,
                 reg62,
                 reg63,
                 reg64,
                 forvar65,
                 reg66,
                 forvar67,
                 reg68,
                 reg69,
                 reg70,
                 reg71,
                 reg72,
                 wire139,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg62 = wire58[(1'h0):(1'h0)];
      reg63 = (wire58[(3'h4):(1'h0)] ?
          {$signed($unsigned(reg62))} : $signed(wire58));
      reg64 <= ({wire60[(3'h4):(2'h2)]} ?
          ((wire58 ?
                  ((wire58 - reg63) ?
                      ((8'hb1) ?
                          reg62 : wire61) : ((8'hb6) ^~ wire59)) : $unsigned((reg63 <<< (7'h44)))) ?
              ({((8'hba) * reg62), {reg63}} ?
                  (wire61 ?
                      $unsigned(wire59) : $signed(wire59)) : wire61) : $unsigned((&$signed(wire58)))) : $unsigned((((|wire59) != reg62[(5'h10):(4'h9)]) < (~|wire60))));
      for (forvar65 = (1'h0); (forvar65 < (1'h0)); forvar65 = (forvar65 + (1'h1)))
        begin
          reg66 <= (&$unsigned({$unsigned($signed(wire60))}));
          for (forvar67 = (1'h0); (forvar67 < (2'h2)); forvar67 = (forvar67 + (1'h1)))
            begin
              reg68 = (^~($signed($signed($unsigned(wire60))) ?
                  wire58 : (^~{$signed(forvar67)})));
            end
          reg69 <= forvar67[(3'h4):(2'h3)];
          reg70 <= {(forvar67[(3'h5):(2'h2)] ?
                  $signed($unsigned((wire60 ?
                      reg66 : reg69))) : reg68[(3'h7):(3'h4)]),
              ((reg64[(4'hb):(4'ha)] ?
                  $signed((reg64 ? reg66 : reg64)) : (~^(wire60 ?
                      wire61 : forvar65))) ^ (8'ha5))};
          reg71 <= (~^($unsigned({$unsigned(reg64)}) ?
              (8'hb1) : $signed($unsigned({wire58, wire58}))));
        end
      reg72 <= reg68[(5'h10):(4'h8)];
    end
  module73 modinst140 (wire139, clk, wire58, reg64, forvar67, reg68, wire60);
  always
    @(posedge clk) begin
      reg141 = (~^$signed(reg64));
      reg142 <= wire59;
      reg143 <= ((^(^~$signed($unsigned((8'hbe))))) ^~ $unsigned(wire61[(2'h2):(1'h1)]));
      reg144 <= $unsigned({((reg64 ?
              $unsigned(reg142) : $signed((8'hb7))) >> ($signed(reg71) ?
              (wire139 << wire59) : (wire59 ? forvar65 : reg142)))});
    end
  assign wire145 = {((8'hbb) && $signed($signed($signed(forvar67))))};
  assign wire146 = reg72[(1'h1):(1'h0)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module73  (y, clk, wire78, wire77, wire76, wire75, wire74);
  output wire [(32'h2ca):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire78;
  input wire [(3'h4):(1'h0)] wire77;
  input wire signed [(4'hd):(1'h0)] wire76;
  input wire signed [(5'h12):(1'h0)] wire75;
  input wire [(4'hc):(1'h0)] wire74;
  wire [(4'ha):(1'h0)] wire138;
  reg signed [(5'h11):(1'h0)] reg137 = (1'h0);
  reg [(4'h8):(1'h0)] reg136 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg135 = (1'h0);
  reg [(4'ha):(1'h0)] reg134 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg133 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar132 = (1'h0);
  reg [(3'h4):(1'h0)] reg131 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire130;
  reg [(4'h8):(1'h0)] reg129 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg128 = (1'h0);
  reg [(5'h12):(1'h0)] reg127 = (1'h0);
  reg [(4'h8):(1'h0)] reg126 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg125 = (1'h0);
  reg [(4'ha):(1'h0)] reg124 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire123;
  reg signed [(5'h15):(1'h0)] reg122 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg121 = (1'h0);
  reg [(4'h9):(1'h0)] reg120 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg119 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg118 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar117 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg116 = (1'h0);
  reg [(4'hf):(1'h0)] reg115 = (1'h0);
  reg [(4'h8):(1'h0)] forvar114 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg113 = (1'h0);
  reg [(2'h3):(1'h0)] reg112 = (1'h0);
  reg [(5'h12):(1'h0)] reg111 = (1'h0);
  reg [(5'h15):(1'h0)] reg110 = (1'h0);
  reg [(5'h10):(1'h0)] forvar109 = (1'h0);
  wire [(5'h14):(1'h0)] wire108;
  reg [(4'hf):(1'h0)] reg107 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar106 = (1'h0);
  reg [(3'h4):(1'h0)] reg105 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire104;
  wire [(3'h6):(1'h0)] wire103;
  reg signed [(3'h4):(1'h0)] reg102 = (1'h0);
  reg [(3'h4):(1'h0)] reg101 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg100 = (1'h0);
  reg [(4'he):(1'h0)] reg99 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg98 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg97 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar96 = (1'h0);
  reg [(3'h5):(1'h0)] reg95 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar94 = (1'h0);
  wire [(5'h12):(1'h0)] wire93;
  reg [(2'h3):(1'h0)] reg92 = (1'h0);
  reg [(3'h4):(1'h0)] reg91 = (1'h0);
  reg [(5'h11):(1'h0)] reg90 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg89 = (1'h0);
  reg [(4'ha):(1'h0)] reg88 = (1'h0);
  reg [(4'hf):(1'h0)] forvar87 = (1'h0);
  reg [(4'hb):(1'h0)] reg86 = (1'h0);
  reg [(5'h12):(1'h0)] reg85 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg84 = (1'h0);
  reg [(3'h5):(1'h0)] forvar83 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg82 = (1'h0);
  reg [(4'hc):(1'h0)] reg81 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg80 = (1'h0);
  wire [(4'ha):(1'h0)] wire79;
  assign y = {wire138,
                 reg137,
                 reg136,
                 reg135,
                 reg134,
                 reg133,
                 forvar132,
                 reg131,
                 wire130,
                 reg129,
                 reg128,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 wire123,
                 reg122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 forvar117,
                 reg116,
                 reg115,
                 forvar114,
                 reg113,
                 reg112,
                 reg111,
                 reg110,
                 forvar109,
                 wire108,
                 reg107,
                 forvar106,
                 reg105,
                 wire104,
                 wire103,
                 reg102,
                 reg101,
                 reg100,
                 reg99,
                 reg98,
                 reg97,
                 forvar96,
                 reg95,
                 forvar94,
                 wire93,
                 reg92,
                 reg91,
                 reg90,
                 reg89,
                 reg88,
                 forvar87,
                 reg86,
                 reg85,
                 reg84,
                 forvar83,
                 reg82,
                 reg81,
                 reg80,
                 wire79,
                 (1'h0)};
  assign wire79 = (~^(wire76 << (&wire77)));
  always
    @(posedge clk) begin
      reg80 = wire76[(3'h5):(2'h3)];
      reg81 <= wire75[(4'hd):(1'h1)];
      reg82 <= ((8'hba) != (8'h9d));
      for (forvar83 = (1'h0); (forvar83 < (2'h2)); forvar83 = (forvar83 + (1'h1)))
        begin
          reg84 <= (((~^wire74[(4'ha):(1'h0)]) ?
                  (reg80 ?
                      forvar83 : $signed(forvar83[(2'h3):(1'h1)])) : {wire75[(3'h4):(3'h4)]}) ?
              (wire79[(3'h5):(1'h0)] + ($signed((forvar83 == wire76)) ?
                  reg80[(3'h7):(1'h1)] : $unsigned((reg80 << wire78)))) : ((^~((8'haa) ~^ (wire78 == wire75))) ?
                  wire78[(1'h1):(1'h1)] : (^(((8'hbc) || wire75) ?
                      reg81[(3'h4):(1'h0)] : $signed(wire78)))));
          reg85 <= {((wire77[(3'h4):(2'h2)] >>> $unsigned(((8'hbd) ?
                      reg84 : wire75))) ?
                  wire79[(3'h4):(1'h1)] : {wire78[(1'h0):(1'h0)],
                      reg82[(1'h0):(1'h0)]}),
              {$signed({(-(8'h9d))}), reg84[(3'h7):(3'h7)]}};
          reg86 <= wire78[(2'h2):(1'h1)];
          for (forvar87 = (1'h0); (forvar87 < (2'h2)); forvar87 = (forvar87 + (1'h1)))
            begin
              reg88 <= $unsigned((^~({$unsigned(wire74),
                  $signed(wire74)} - $signed(reg84))));
              reg89 <= (~^{wire78[(3'h6):(1'h1)],
                  $unsigned($signed($signed(wire77)))});
              reg90 <= $signed($signed($unsigned(wire78[(3'h4):(1'h1)])));
            end
          reg91 = (+wire76[(3'h5):(1'h0)]);
        end
    end
  always
    @(posedge clk) begin
      reg92 = (~|(8'hac));
    end
  assign wire93 = reg82;
  always
    @(posedge clk) begin
      for (forvar94 = (1'h0); (forvar94 < (1'h1)); forvar94 = (forvar94 + (1'h1)))
        begin
          reg95 = {reg89,
              (+(((8'hb1) ? (~&reg92) : forvar83[(1'h0):(1'h0)]) ?
                  wire93[(2'h3):(2'h3)] : {$signed(reg89), reg89}))};
          for (forvar96 = (1'h0); (forvar96 < (2'h2)); forvar96 = (forvar96 + (1'h1)))
            begin
              reg97 <= forvar94[(2'h3):(2'h2)];
              reg98 <= (reg92 >> ($unsigned($unsigned((wire93 ?
                  forvar87 : wire76))) <<< forvar96[(5'h10):(4'ha)]));
              reg99 <= (^~reg88);
              reg100 <= wire78[(4'h8):(2'h2)];
            end
          reg101 <= {((&$unsigned($unsigned(reg82))) <= wire93),
              $unsigned($unsigned(reg84))};
          reg102 <= reg99[(4'he):(2'h2)];
        end
    end
  assign wire103 = reg99;
  assign wire104 = $signed((reg102 ?
                       $unsigned(((reg89 && (8'hb5)) ?
                           forvar96 : forvar94)) : reg101[(3'h4):(2'h3)]));
  always
    @(posedge clk) begin
      reg105 <= (&$signed($unsigned(($unsigned(wire74) ?
          (wire79 ? reg98 : reg100) : $signed(forvar94)))));
      for (forvar106 = (1'h0); (forvar106 < (1'h0)); forvar106 = (forvar106 + (1'h1)))
        begin
          reg107 = {(reg105 ?
                  $signed(reg88[(3'h5):(3'h4)]) : reg86[(4'hb):(4'hb)])};
        end
    end
  assign wire108 = {$unsigned($signed($unsigned((reg100 ? reg80 : reg100)))),
                       (^wire75[(3'h7):(3'h7)])};
  always
    @(posedge clk) begin
      for (forvar109 = (1'h0); (forvar109 < (2'h2)); forvar109 = (forvar109 + (1'h1)))
        begin
          reg110 = ((wire103 >= (~&$unsigned($signed((8'ha1))))) ?
              $unsigned($signed(((reg98 ? wire77 : reg85) ?
                  (reg101 ?
                      forvar87 : reg81) : forvar109))) : $unsigned(((reg80[(3'h5):(3'h4)] != reg88) ?
                  reg91 : $signed($signed(wire104)))));
          reg111 = wire103[(2'h2):(1'h0)];
          reg112 <= $unsigned({$signed($signed((reg81 ? reg101 : forvar87))),
              (wire104 ?
                  (wire75[(3'h7):(1'h1)] ?
                      $unsigned(wire77) : (reg99 & wire103)) : (&$unsigned((8'hbe))))});
        end
      reg113 = ($signed((reg100 ?
          $unsigned($unsigned(reg99)) : $unsigned((&reg102)))) >> (($signed({(8'h9d),
          forvar106}) & wire77) ~^ $unsigned($unsigned({forvar83, forvar87}))));
      for (forvar114 = (1'h0); (forvar114 < (1'h1)); forvar114 = (forvar114 + (1'h1)))
        begin
          reg115 = forvar114[(3'h5):(1'h1)];
          reg116 <= $unsigned({((^{wire79, forvar87}) ?
                  (reg97[(1'h1):(1'h1)] ?
                      (reg86 ?
                          wire104 : reg115) : (8'hb7)) : $signed(reg99[(4'hd):(3'h7)])),
              (|((~|reg110) ? $unsigned(reg90) : (reg80 * reg92)))});
        end
    end
  always
    @(posedge clk) begin
      for (forvar117 = (1'h0); (forvar117 < (2'h3)); forvar117 = (forvar117 + (1'h1)))
        begin
          reg118 = reg101;
          reg119 <= wire103[(3'h5):(1'h0)];
          reg120 <= $unsigned($unsigned(($signed($signed((8'had))) ?
              $unsigned((wire76 ?
                  (8'hb9) : forvar94)) : (~|(wire108 & (8'hb5))))));
          reg121 <= (~$unsigned(forvar83[(1'h1):(1'h1)]));
        end
      reg122 <= (-{(forvar114 ?
              reg105[(2'h3):(1'h1)] : (forvar94[(3'h7):(3'h4)] ?
                  {reg111} : $signed(wire75)))});
    end
  assign wire123 = (reg120[(2'h2):(1'h0)] ?
                       $unsigned(wire79[(3'h5):(2'h3)]) : forvar106[(2'h3):(2'h3)]);
  always
    @(posedge clk) begin
      reg124 <= (~(forvar106 ?
          $unsigned({((8'hb1) ? reg111 : reg100)}) : reg111));
      reg125 <= ((-$signed(reg101)) ? reg115 : forvar117);
      reg126 <= reg89;
      reg127 <= (~^($unsigned($signed(wire75[(1'h1):(1'h1)])) ?
          (((wire74 ? reg89 : reg84) >>> (reg97 ?
              reg88 : (8'ha4))) - reg97[(1'h1):(1'h1)]) : wire108));
    end
  always
    @(posedge clk) begin
      reg128 <= {wire93, wire77};
      reg129 = $unsigned($signed($unsigned(($signed(reg124) - $signed(reg86)))));
    end
  assign wire130 = (reg102 ?
                       (reg102[(1'h1):(1'h0)] ?
                           {$signed((reg80 == reg95)),
                               (&((7'h43) ?
                                   reg110 : reg90))} : {{(reg119 <= reg125),
                                   $signed(forvar117)}}) : (^wire104[(3'h5):(3'h4)]));
  always
    @(posedge clk) begin
      reg131 <= $signed((+$signed(((reg110 ? reg98 : wire77) ?
          $unsigned(reg101) : reg116))));
      for (forvar132 = (1'h0); (forvar132 < (2'h3)); forvar132 = (forvar132 + (1'h1)))
        begin
          reg133 <= (-$signed($unsigned($unsigned((~^reg105)))));
        end
      reg134 <= $signed($unsigned((((reg110 & (8'hb8)) && $unsigned((8'hb5))) | ($unsigned(reg119) >= (~^wire79)))));
      reg135 <= reg110[(1'h0):(1'h0)];
      reg136 <= $unsigned(((~(8'ha2)) | (+(((8'ha2) < reg112) > (forvar83 <= (8'ha3))))));
    end
  always
    @(posedge clk) begin
      reg137 <= $signed(($signed(($signed((8'ha2)) ?
          {reg98} : $signed(wire77))) >= $signed(($signed(reg129) ^~ (reg122 ?
          reg112 : (7'h40))))));
    end
  assign wire138 = ({(reg127[(3'h6):(3'h5)] <<< wire77[(1'h1):(1'h1)])} * reg134[(3'h4):(1'h1)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module213
#( parameter param459 = (((~&(!{(7'h41)})) != ((~&(!(8'ha8))) <<< {((8'had) ? (7'h44) : (8'ha2))})) - (!(!((~|(8'hb1)) >= (~^(8'had)))))) )
(y, clk, wire217, wire216, wire215, wire214);
  output wire [(32'h1d3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire217;
  input wire signed [(5'h11):(1'h0)] wire216;
  input wire signed [(2'h2):(1'h0)] wire215;
  input wire signed [(2'h3):(1'h0)] wire214;
  reg [(4'he):(1'h0)] reg458 = (1'h0);
  reg [(3'h5):(1'h0)] reg457 = (1'h0);
  reg [(4'h9):(1'h0)] reg456 = (1'h0);
  reg [(5'h12):(1'h0)] reg455 = (1'h0);
  reg [(4'hf):(1'h0)] reg454 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg453 = (1'h0);
  reg [(3'h4):(1'h0)] reg452 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg451 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg450 = (1'h0);
  wire [(4'h8):(1'h0)] wire449;
  wire [(5'h11):(1'h0)] wire448;
  wire signed [(4'hd):(1'h0)] wire349;
  wire [(5'h14):(1'h0)] wire231;
  reg signed [(4'hf):(1'h0)] reg230 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg229 = (1'h0);
  reg [(4'he):(1'h0)] reg228 = (1'h0);
  reg [(5'h12):(1'h0)] reg227 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg226 = (1'h0);
  reg [(4'h9):(1'h0)] forvar225 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg224 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg223 = (1'h0);
  reg [(4'hf):(1'h0)] reg222 = (1'h0);
  reg [(4'he):(1'h0)] reg221 = (1'h0);
  reg [(5'h15):(1'h0)] reg220 = (1'h0);
  reg [(5'h14):(1'h0)] forvar219 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg218 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire351;
  reg signed [(4'h9):(1'h0)] reg352 = (1'h0);
  reg [(4'he):(1'h0)] reg353 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg354 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg355 = (1'h0);
  reg signed [(4'he):(1'h0)] reg356 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg357 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg358 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg359 = (1'h0);
  reg [(5'h14):(1'h0)] reg360 = (1'h0);
  reg [(3'h4):(1'h0)] reg361 = (1'h0);
  reg [(3'h4):(1'h0)] reg362 = (1'h0);
  wire [(2'h3):(1'h0)] wire446;
  assign y = {reg458,
                 reg457,
                 reg456,
                 reg455,
                 reg454,
                 reg453,
                 reg452,
                 reg451,
                 reg450,
                 wire449,
                 wire448,
                 wire349,
                 wire231,
                 reg230,
                 reg229,
                 reg228,
                 reg227,
                 reg226,
                 forvar225,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 forvar219,
                 reg218,
                 wire351,
                 reg352,
                 reg353,
                 reg354,
                 reg355,
                 reg356,
                 reg357,
                 reg358,
                 reg359,
                 reg360,
                 reg361,
                 reg362,
                 wire446,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg218 <= wire217[(2'h3):(1'h1)];
      for (forvar219 = (1'h0); (forvar219 < (1'h1)); forvar219 = (forvar219 + (1'h1)))
        begin
          reg220 = $signed((wire214[(2'h3):(2'h2)] ~^ ({(8'ha0),
                  $unsigned(reg218)} ?
              (-$signed(forvar219)) : (|{wire216, forvar219}))));
          reg221 = (reg220 | ($signed(wire216) <<< $signed($unsigned(forvar219[(1'h0):(1'h0)]))));
          reg222 <= wire217;
          reg223 <= $signed($signed((|reg221)));
          reg224 = {wire214[(1'h1):(1'h1)], (8'hae)};
        end
      for (forvar225 = (1'h0); (forvar225 < (1'h1)); forvar225 = (forvar225 + (1'h1)))
        begin
          reg226 <= reg218[(2'h2):(1'h0)];
          reg227 <= (8'hba);
          reg228 <= wire214;
        end
      reg229 <= (8'hb3);
      reg230 <= {(7'h42)};
    end
  assign wire231 = (forvar219[(3'h5):(3'h4)] ?
                       (wire215 == reg230) : $unsigned(($signed((reg227 ?
                           reg230 : wire217)) << (wire214 ~^ $unsigned(wire216)))));
  module232 modinst350 (wire349, clk, wire217, wire216, reg221, forvar219, reg228);
  assign wire351 = $unsigned(((^forvar225[(1'h1):(1'h0)]) ?
                       $signed({(~|reg226)}) : (($signed(wire217) * reg223) - $unsigned($unsigned(wire214)))));
  always
    @(posedge clk) begin
      reg352 = $signed({($signed((forvar225 ?
              reg223 : (8'hb2))) ^~ $unsigned((wire214 ? reg230 : reg226)))});
      reg353 <= {$signed(reg218)};
    end
  always
    @(posedge clk) begin
      reg354 <= $signed($unsigned(($signed((!(8'ha2))) ?
          wire216[(3'h6):(3'h5)] : reg229[(1'h0):(1'h0)])));
      reg355 <= reg230[(4'h9):(4'h9)];
      reg356 <= {$signed((8'had))};
      reg357 = ((reg355[(2'h2):(1'h0)] > $signed((^~reg223[(3'h5):(3'h5)]))) >= (~({(~|reg226),
          (reg355 ? wire214 : reg355)} || forvar219)));
      reg358 = reg357;
    end
  always
    @(posedge clk) begin
      reg359 <= $unsigned((((8'hb2) ^ $unsigned((~|reg221))) ?
          ($signed($signed(reg354)) <= $signed(wire349[(2'h2):(2'h2)])) : reg227[(2'h3):(2'h2)]));
    end
  always
    @(posedge clk) begin
      reg360 <= wire214;
      reg361 <= (reg356[(3'h5):(2'h3)] ?
          ({reg223} ?
              reg230[(4'h8):(3'h4)] : reg358[(3'h6):(2'h2)]) : (+($unsigned(reg353) <<< ((8'ha2) ?
              (reg356 != (8'hb2)) : (reg357 ? reg228 : reg221)))));
      reg362 <= (|$unsigned((&(~&(~|reg356)))));
    end
  module363 modinst447 (wire446, clk, wire217, wire231, reg224, reg357, reg358);
  assign wire448 = ({(~((reg359 ? reg355 : reg223) ? {wire446} : (^reg353))),
                           $unsigned(($unsigned(reg354) <<< wire215[(2'h2):(2'h2)]))} ?
                       $unsigned((^forvar219)) : ($unsigned(wire215) + $unsigned(($signed(reg229) ?
                           (reg226 ?
                               wire215 : reg222) : reg362[(3'h4):(1'h0)]))));
  assign wire449 = $unsigned(reg220[(4'hc):(3'h7)]);
  always
    @(posedge clk) begin
      if (wire214)
        begin
          reg450 = ((reg227[(5'h10):(1'h1)] | reg356) ?
              ($signed(reg356) - (+(^~(+wire351)))) : ($signed((^(wire349 ~^ reg224))) <<< ($unsigned($signed(reg357)) == (-reg360[(1'h1):(1'h1)]))));
        end
      else
        begin
          reg450 <= (-($signed((~$unsigned(wire217))) | ((-((8'hb3) >= (8'ha6))) - ($unsigned(reg359) ?
              {wire216, (8'h9d)} : (wire448 + reg450)))));
          reg451 <= reg360;
          reg452 <= ((wire214[(2'h3):(1'h0)] || reg221) ?
              forvar225[(2'h3):(2'h3)] : $unsigned(((~&reg352) & $unsigned((reg362 << reg355)))));
          reg453 <= $unsigned((reg451[(3'h6):(2'h2)] - $signed((+$unsigned(reg221)))));
        end
    end
  always
    @(posedge clk) begin
      reg454 <= $signed($unsigned(forvar219));
      reg455 <= ((!($signed($signed(reg357)) * (~|reg230[(4'he):(4'ha)]))) && reg450[(1'h1):(1'h0)]);
      reg456 <= (^~($signed({(reg221 ? (8'ha3) : reg453),
              reg360[(5'h12):(4'hf)]}) ?
          (~^$signed(reg452)) : (($signed(wire349) ?
              {reg218} : {(8'haf)}) != reg353[(3'h6):(1'h0)])));
      reg457 <= (reg222[(2'h2):(1'h0)] ?
          {(wire448[(5'h10):(2'h3)] ?
                  (reg356 ~^ (wire217 ? (8'hb0) : reg354)) : $signed({reg356,
                      reg359}))} : $unsigned(wire231[(4'h9):(4'h8)]));
      reg458 <= reg230[(3'h5):(1'h1)];
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module363
#( parameter param444 = {(&(((8'h9c) == ((8'hac) ? (8'hbc) : (8'ha5))) ? (|((8'ha4) ? (8'hab) : (8'h9e))) : {{(7'h40)}, ((8'hb7) ? (8'ha8) : (8'hb6))}))}
, parameter param445 = ((~param444) ? param444 : (({(param444 ? param444 : param444), (param444 ? (8'h9d) : param444)} | (param444 ? (param444 + param444) : (param444 ? param444 : param444))) >>> (((+param444) > {param444}) == (&((8'ha1) ? param444 : param444))))) )
(y, clk, wire368, wire367, wire366, wire365, wire364);
  output wire [(32'h341):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire368;
  input wire [(5'h13):(1'h0)] wire367;
  input wire signed [(4'ha):(1'h0)] wire366;
  input wire [(2'h3):(1'h0)] wire365;
  input wire signed [(2'h3):(1'h0)] wire364;
  reg signed [(5'h13):(1'h0)] reg443 = (1'h0);
  reg [(3'h7):(1'h0)] reg442 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg441 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg440 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar439 = (1'h0);
  reg [(4'hc):(1'h0)] reg438 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg437 = (1'h0);
  reg [(3'h7):(1'h0)] reg436 = (1'h0);
  reg [(4'hb):(1'h0)] reg435 = (1'h0);
  reg [(2'h2):(1'h0)] reg434 = (1'h0);
  reg [(2'h2):(1'h0)] forvar433 = (1'h0);
  wire [(4'ha):(1'h0)] wire432;
  wire [(5'h10):(1'h0)] wire431;
  wire [(4'hf):(1'h0)] wire430;
  reg [(5'h15):(1'h0)] reg429 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg428 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg427 = (1'h0);
  reg [(3'h4):(1'h0)] reg426 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg425 = (1'h0);
  reg [(3'h5):(1'h0)] reg424 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar423 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar422 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg421 = (1'h0);
  reg [(5'h14):(1'h0)] reg420 = (1'h0);
  reg [(4'he):(1'h0)] reg419 = (1'h0);
  reg [(5'h12):(1'h0)] reg418 = (1'h0);
  wire [(4'hf):(1'h0)] wire417;
  wire [(5'h12):(1'h0)] wire416;
  wire signed [(3'h5):(1'h0)] wire415;
  reg [(4'hb):(1'h0)] reg414 = (1'h0);
  reg [(3'h7):(1'h0)] reg413 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg412 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar411 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg410 = (1'h0);
  reg [(4'hc):(1'h0)] reg409 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg408 = (1'h0);
  reg [(5'h11):(1'h0)] reg407 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg406 = (1'h0);
  reg [(4'hb):(1'h0)] reg405 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar404 = (1'h0);
  reg [(4'h9):(1'h0)] reg403 = (1'h0);
  reg [(4'hd):(1'h0)] reg402 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg401 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg400 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg399 = (1'h0);
  reg [(5'h15):(1'h0)] reg398 = (1'h0);
  reg [(3'h4):(1'h0)] reg397 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar396 = (1'h0);
  reg [(4'he):(1'h0)] reg395 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg394 = (1'h0);
  wire [(4'ha):(1'h0)] wire393;
  reg [(4'hb):(1'h0)] reg392 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar391 = (1'h0);
  reg [(5'h15):(1'h0)] reg390 = (1'h0);
  reg [(5'h13):(1'h0)] reg389 = (1'h0);
  reg [(5'h15):(1'h0)] reg388 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg387 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg386 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg385 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire384;
  reg [(3'h5):(1'h0)] reg383 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg382 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg381 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg380 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar379 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg378 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg377 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar376 = (1'h0);
  reg [(2'h3):(1'h0)] reg375 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg374 = (1'h0);
  wire [(3'h5):(1'h0)] wire373;
  reg signed [(3'h4):(1'h0)] reg372 = (1'h0);
  reg [(5'h15):(1'h0)] reg371 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg370 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg369 = (1'h0);
  assign y = {reg443,
                 reg442,
                 reg441,
                 reg440,
                 forvar439,
                 reg438,
                 reg437,
                 reg436,
                 reg435,
                 reg434,
                 forvar433,
                 wire432,
                 wire431,
                 wire430,
                 reg429,
                 reg428,
                 reg427,
                 reg426,
                 reg425,
                 reg424,
                 forvar423,
                 forvar422,
                 reg421,
                 reg420,
                 reg419,
                 reg418,
                 wire417,
                 wire416,
                 wire415,
                 reg414,
                 reg413,
                 reg412,
                 forvar411,
                 reg410,
                 reg409,
                 reg408,
                 reg407,
                 reg406,
                 reg405,
                 forvar404,
                 reg403,
                 reg402,
                 reg401,
                 reg400,
                 reg399,
                 reg398,
                 reg397,
                 forvar396,
                 reg395,
                 reg394,
                 wire393,
                 reg392,
                 forvar391,
                 reg390,
                 reg389,
                 reg388,
                 reg387,
                 reg386,
                 reg385,
                 wire384,
                 reg383,
                 reg382,
                 reg381,
                 reg380,
                 forvar379,
                 reg378,
                 reg377,
                 forvar376,
                 reg375,
                 reg374,
                 wire373,
                 reg372,
                 reg371,
                 reg370,
                 reg369,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg369 <= (8'hb9);
      reg370 = $unsigned($unsigned($signed((-$unsigned(wire364)))));
      reg371 = (~&{(($signed(wire364) ?
                  wire367[(4'he):(4'ha)] : wire368[(2'h3):(1'h1)]) ?
              (8'hb3) : (wire364 ?
                  ((8'hb3) ? reg370 : (8'had)) : (wire367 << wire366))),
          reg370[(4'h8):(2'h3)]});
      reg372 <= (-(~|$unsigned((^~(~^wire366)))));
    end
  assign wire373 = reg372[(2'h2):(1'h0)];
  always
    @(posedge clk) begin
      reg374 <= $unsigned(wire368);
      reg375 <= wire365;
      for (forvar376 = (1'h0); (forvar376 < (2'h3)); forvar376 = (forvar376 + (1'h1)))
        begin
          reg377 = (-wire373[(1'h0):(1'h0)]);
          reg378 <= ($signed($signed({$unsigned(reg374),
              reg369})) || $unsigned((|($unsigned((8'ha0)) <= (&wire365)))));
          for (forvar379 = (1'h0); (forvar379 < (3'h4)); forvar379 = (forvar379 + (1'h1)))
            begin
              reg380 <= wire368[(1'h1):(1'h1)];
              reg381 <= $unsigned($signed((wire368 - $signed((reg380 ^ forvar379)))));
            end
          reg382 <= (~&{$unsigned({forvar376, $unsigned((8'h9f))}), wire368});
          reg383 <= $signed(reg371);
        end
    end
  assign wire384 = $signed($unsigned(forvar379[(4'hb):(1'h1)]));
  always
    @(posedge clk) begin
      reg385 <= reg370;
      reg386 <= ((~($unsigned((reg371 ~^ reg369)) ?
          $unsigned(wire373[(1'h0):(1'h0)]) : wire367)) >>> {$unsigned(((reg374 <<< wire364) >= (reg377 ?
              wire373 : reg381))),
          forvar376[(3'h5):(1'h0)]});
      reg387 <= reg382[(3'h5):(1'h1)];
      reg388 <= (-{(&$signed($signed((8'ha1))))});
      reg389 = wire368[(3'h5):(3'h5)];
    end
  always
    @(posedge clk) begin
      reg390 = $unsigned((~^reg382));
      for (forvar391 = (1'h0); (forvar391 < (2'h3)); forvar391 = (forvar391 + (1'h1)))
        begin
          reg392 <= reg386[(4'hb):(1'h0)];
        end
    end
  assign wire393 = ((8'haf) ?
                       (&$signed($signed((~^reg386)))) : reg383[(1'h1):(1'h1)]);
  always
    @(posedge clk) begin
      reg394 <= wire364[(2'h2):(2'h2)];
      reg395 <= $unsigned((~&reg394[(1'h1):(1'h0)]));
      for (forvar396 = (1'h0); (forvar396 < (3'h4)); forvar396 = (forvar396 + (1'h1)))
        begin
          reg397 <= $unsigned(($unsigned(reg378) <<< (reg377[(4'hf):(3'h6)] ?
              $signed({reg375, reg383}) : wire367)));
          if (($unsigned(wire367) >>> $unsigned($unsigned($signed($signed(wire365))))))
            begin
              reg398 = $unsigned(reg369);
              reg399 = {$signed({$signed((-wire368)),
                      (reg371 ? $unsigned(reg370) : ((8'hba) != reg369))}),
                  ({($signed(wire366) ? reg387 : $signed(forvar396)),
                      reg397[(3'h4):(2'h3)]} <= {(+(wire365 || (8'hbd)))})};
              reg400 = $signed(reg371[(4'hb):(4'h8)]);
              reg401 <= {((8'hae) != ((~reg374[(3'h7):(1'h1)]) ?
                      (wire384 ?
                          reg388 : $signed(wire365)) : $signed($unsigned(reg398))))};
              reg402 = $signed($unsigned((^~reg397)));
            end
          else
            begin
              reg398 <= forvar379;
            end
          reg403 <= $unsigned((reg401[(3'h7):(2'h3)] ~^ (wire366 ?
              (-$unsigned(reg377)) : (reg370[(2'h3):(2'h3)] ?
                  wire366 : $signed(reg389)))));
        end
      for (forvar404 = (1'h0); (forvar404 < (3'h4)); forvar404 = (forvar404 + (1'h1)))
        begin
          reg405 = $unsigned(((((|forvar404) ?
                  $unsigned(reg399) : (~reg372)) >> ((+reg387) ?
                  ((8'hb3) ? wire364 : reg378) : (wire384 ?
                      reg372 : forvar404))) ?
              $unsigned(forvar404) : reg386));
        end
    end
  always
    @(posedge clk) begin
      reg406 <= (8'hb3);
      reg407 = (&(reg400[(1'h1):(1'h1)] - $unsigned(($unsigned(reg395) ?
          (wire368 > forvar391) : $signed(reg402)))));
      reg408 = forvar396[(2'h2):(2'h2)];
      reg409 <= forvar379;
      reg410 <= (&(8'hbe));
    end
  always
    @(posedge clk) begin
      for (forvar411 = (1'h0); (forvar411 < (1'h1)); forvar411 = (forvar411 + (1'h1)))
        begin
          reg412 = $unsigned($unsigned((((!wire365) ?
              (reg374 ?
                  reg409 : reg406) : (~^reg370)) * (&reg383[(3'h5):(3'h4)]))));
        end
      reg413 <= ($unsigned($signed(reg410)) ?
          reg388[(3'h6):(3'h6)] : {(~&{(!(8'h9f))}),
              (((!(8'ha8)) != $unsigned((8'hb5))) || forvar376)});
      reg414 <= reg405[(2'h3):(2'h3)];
    end
  assign wire415 = $unsigned(forvar404);
  assign wire416 = wire415;
  assign wire417 = $unsigned((~|$signed(reg401[(4'ha):(2'h2)])));
  always
    @(posedge clk) begin
      reg418 <= (-((+($signed(reg392) ?
          (|wire393) : {wire415, reg375})) + (+wire367)));
      reg419 = (($unsigned($unsigned((reg370 ? reg374 : reg380))) != reg394) ?
          reg387[(4'ha):(1'h1)] : $unsigned((~&$unsigned($signed(wire415)))));
      reg420 <= $signed((forvar404[(3'h5):(2'h3)] ?
          $signed(forvar404[(2'h2):(1'h1)]) : $unsigned((+reg371))));
      reg421 <= (~^(^$unsigned({(reg413 ? forvar411 : reg372)})));
    end
  always
    @(posedge clk) begin
      for (forvar422 = (1'h0); (forvar422 < (1'h1)); forvar422 = (forvar422 + (1'h1)))
        begin
          for (forvar423 = (1'h0); (forvar423 < (3'h4)); forvar423 = (forvar423 + (1'h1)))
            begin
              reg424 <= $signed(reg413);
            end
          reg425 = ($signed(($signed({reg398}) << reg418)) ^~ $unsigned((wire415[(1'h0):(1'h0)] > reg401[(1'h1):(1'h0)])));
        end
      reg426 <= wire366;
      reg427 <= (&((reg419 << (reg387 ?
          reg394 : (~^forvar404))) - wire364[(1'h0):(1'h0)]));
      reg428 <= forvar422[(1'h0):(1'h0)];
      reg429 <= (forvar404 & {(reg390[(3'h5):(2'h2)] || $unsigned((forvar391 ?
              (8'hbf) : reg387))),
          reg394});
    end
  assign wire430 = ($signed(((+(reg371 ^ reg377)) ?
                       ((reg421 ? wire366 : forvar391) ?
                           reg386 : (!(8'ha2))) : reg395)) & (((-{(8'h9f)}) ?
                       $signed(reg429[(1'h0):(1'h0)]) : $signed((reg383 >>> forvar422))) ^~ (^~forvar411[(3'h5):(1'h0)])));
  assign wire431 = ((reg405[(4'h8):(2'h3)] ?
                           (reg406[(2'h3):(1'h1)] <= (~&((8'hb3) ?
                               forvar404 : wire415))) : wire368[(1'h0):(1'h0)]) ?
                       $unsigned((reg374 ?
                           forvar411[(1'h1):(1'h0)] : {(-reg394),
                               ((8'h9e) ? forvar376 : reg428)})) : (reg372 ?
                           $signed($signed((~&reg401))) : (&(wire373 | (~^forvar411)))));
  assign wire432 = (wire393 ?
                       ((reg380[(4'hd):(4'h8)] ?
                           $signed(wire367[(3'h6):(1'h1)]) : ({reg410} & reg387)) || reg429) : (8'hb0));
  always
    @(posedge clk) begin
      for (forvar433 = (1'h0); (forvar433 < (1'h0)); forvar433 = (forvar433 + (1'h1)))
        begin
          reg434 <= ($signed({$signed({wire365}),
              reg382}) ^ forvar404[(2'h3):(1'h0)]);
          reg435 = ($signed(((wire393 ?
              wire373[(1'h0):(1'h0)] : (forvar379 > reg401)) > (wire393 ?
              $signed(reg434) : {reg429, reg403}))) && reg374);
          reg436 = $signed(reg378[(2'h3):(1'h0)]);
          reg437 <= ((^~($signed({reg369, wire416}) ?
                  $signed($unsigned((8'hb2))) : (-(forvar433 != reg428)))) ?
              (($signed((reg370 ? (7'h40) : reg434)) ?
                      ((reg400 ? reg372 : wire368) ?
                          (reg378 != forvar411) : {reg426}) : $unsigned(reg410[(3'h6):(3'h6)])) ?
                  (8'hbb) : forvar404) : $signed(reg377));
          reg438 <= reg392[(1'h1):(1'h0)];
        end
      for (forvar439 = (1'h0); (forvar439 < (1'h1)); forvar439 = (forvar439 + (1'h1)))
        begin
          reg440 <= ((-({reg438[(3'h7):(1'h0)]} == ((reg435 << wire384) ?
              ((8'ha3) ?
                  forvar439 : reg399) : $signed(wire364)))) != $signed($signed({{(8'h9d),
                  forvar391}})));
          reg441 <= reg378;
          reg442 <= {$signed({(8'h9f)})};
          reg443 <= $signed({forvar404[(2'h2):(1'h0)]});
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module232
#( parameter param347 = {((({(7'h44), (8'ha7)} ? (^~(8'ha4)) : (8'hb6)) >> {((7'h43) && (7'h43))}) ? ((!((8'ha7) ? (8'hb0) : (8'ha5))) ^~ ((-(8'hac)) ? ((8'hb9) | (8'had)) : ((8'ha8) ? (8'hb0) : (8'hb5)))) : {{((8'hb3) ? (8'ha0) : (7'h41))}, (7'h42)})}
, parameter param348 = param347 )
(y, clk, wire237, wire236, wire235, wire234, wire233);
  output wire [(32'h4da):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire237;
  input wire signed [(2'h3):(1'h0)] wire236;
  input wire signed [(4'he):(1'h0)] wire235;
  input wire signed [(5'h14):(1'h0)] wire234;
  input wire signed [(4'h8):(1'h0)] wire233;
  reg signed [(5'h15):(1'h0)] reg346 = (1'h0);
  reg [(2'h3):(1'h0)] reg345 = (1'h0);
  reg [(2'h2):(1'h0)] reg344 = (1'h0);
  reg [(4'hf):(1'h0)] reg343 = (1'h0);
  reg [(2'h2):(1'h0)] forvar342 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg341 = (1'h0);
  reg [(2'h2):(1'h0)] reg340 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg339 = (1'h0);
  reg [(5'h15):(1'h0)] reg338 = (1'h0);
  reg [(4'hc):(1'h0)] reg337 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg336 = (1'h0);
  reg [(5'h15):(1'h0)] reg335 = (1'h0);
  reg [(4'hf):(1'h0)] reg334 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg333 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg332 = (1'h0);
  reg [(3'h5):(1'h0)] reg331 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg330 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg329 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg328 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg327 = (1'h0);
  reg [(4'hb):(1'h0)] reg326 = (1'h0);
  reg [(2'h3):(1'h0)] forvar325 = (1'h0);
  reg [(4'he):(1'h0)] reg324 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg323 = (1'h0);
  reg [(4'hd):(1'h0)] reg322 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar321 = (1'h0);
  reg [(4'ha):(1'h0)] reg320 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg319 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg318 = (1'h0);
  reg [(5'h12):(1'h0)] reg317 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg316 = (1'h0);
  reg [(5'h14):(1'h0)] reg315 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg314 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar313 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire312;
  reg [(5'h14):(1'h0)] reg311 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg310 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire309;
  reg [(4'ha):(1'h0)] reg308 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg307 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg306 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg305 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg304 = (1'h0);
  reg [(5'h15):(1'h0)] reg303 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg302 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg301 = (1'h0);
  reg [(5'h14):(1'h0)] reg300 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar299 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire298;
  reg [(5'h10):(1'h0)] reg297 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg296 = (1'h0);
  reg [(4'h9):(1'h0)] reg295 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar294 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg293 = (1'h0);
  reg [(5'h15):(1'h0)] reg292 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg291 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg290 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar289 = (1'h0);
  reg [(5'h13):(1'h0)] reg288 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg287 = (1'h0);
  reg [(5'h12):(1'h0)] reg286 = (1'h0);
  reg [(4'he):(1'h0)] reg285 = (1'h0);
  reg [(4'hf):(1'h0)] reg284 = (1'h0);
  reg [(4'hb):(1'h0)] forvar283 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg282 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg281 = (1'h0);
  reg [(3'h4):(1'h0)] reg280 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg279 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg278 = (1'h0);
  reg [(3'h5):(1'h0)] reg277 = (1'h0);
  reg signed [(4'he):(1'h0)] reg276 = (1'h0);
  reg [(3'h6):(1'h0)] reg275 = (1'h0);
  reg [(4'h9):(1'h0)] reg274 = (1'h0);
  reg [(5'h10):(1'h0)] forvar273 = (1'h0);
  reg signed [(4'he):(1'h0)] reg272 = (1'h0);
  reg [(4'hd):(1'h0)] reg271 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg270 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg269 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar268 = (1'h0);
  reg [(5'h10):(1'h0)] forvar267 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg266 = (1'h0);
  reg [(3'h7):(1'h0)] reg265 = (1'h0);
  reg [(3'h5):(1'h0)] reg264 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg263 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg262 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg261 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg260 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire259;
  reg signed [(4'h9):(1'h0)] reg258 = (1'h0);
  reg [(4'hf):(1'h0)] reg257 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg256 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg255 = (1'h0);
  reg [(3'h6):(1'h0)] reg254 = (1'h0);
  reg [(4'h8):(1'h0)] reg253 = (1'h0);
  reg [(4'h8):(1'h0)] forvar252 = (1'h0);
  reg [(4'hc):(1'h0)] reg251 = (1'h0);
  reg [(4'h8):(1'h0)] forvar250 = (1'h0);
  reg [(4'hf):(1'h0)] reg249 = (1'h0);
  reg [(4'ha):(1'h0)] reg248 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire247;
  reg signed [(5'h11):(1'h0)] reg246 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg245 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar244 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg243 = (1'h0);
  reg [(3'h6):(1'h0)] reg242 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg241 = (1'h0);
  reg [(5'h13):(1'h0)] reg240 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg239 = (1'h0);
  reg [(3'h7):(1'h0)] reg238 = (1'h0);
  assign y = {reg346,
                 reg345,
                 reg344,
                 reg343,
                 forvar342,
                 reg341,
                 reg340,
                 reg339,
                 reg338,
                 reg337,
                 reg336,
                 reg335,
                 reg334,
                 reg333,
                 reg332,
                 reg331,
                 reg330,
                 reg329,
                 reg328,
                 reg327,
                 reg326,
                 forvar325,
                 reg324,
                 reg323,
                 reg322,
                 forvar321,
                 reg320,
                 reg319,
                 reg318,
                 reg317,
                 reg316,
                 reg315,
                 reg314,
                 forvar313,
                 wire312,
                 reg311,
                 reg310,
                 wire309,
                 reg308,
                 reg307,
                 reg306,
                 reg305,
                 reg304,
                 reg303,
                 reg302,
                 reg301,
                 reg300,
                 forvar299,
                 wire298,
                 reg297,
                 reg296,
                 reg295,
                 forvar294,
                 reg293,
                 reg292,
                 reg291,
                 reg290,
                 forvar289,
                 reg288,
                 reg287,
                 reg286,
                 reg285,
                 reg284,
                 forvar283,
                 reg282,
                 reg281,
                 reg280,
                 reg279,
                 reg278,
                 reg277,
                 reg276,
                 reg275,
                 reg274,
                 forvar273,
                 reg272,
                 reg271,
                 reg270,
                 reg269,
                 forvar268,
                 forvar267,
                 reg266,
                 reg265,
                 reg264,
                 reg263,
                 reg262,
                 reg261,
                 reg260,
                 wire259,
                 reg258,
                 reg257,
                 reg256,
                 reg255,
                 reg254,
                 reg253,
                 forvar252,
                 reg251,
                 forvar250,
                 reg249,
                 reg248,
                 wire247,
                 reg246,
                 reg245,
                 forvar244,
                 reg243,
                 reg242,
                 reg241,
                 reg240,
                 reg239,
                 reg238,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg238 <= wire237;
      reg239 <= wire237[(4'ha):(2'h2)];
      reg240 = $unsigned((&(^~$signed((+reg238)))));
      reg241 <= (((8'ha5) ?
          (({reg239, reg240} ?
              $unsigned(reg240) : reg240[(2'h2):(1'h0)]) < wire237) : reg240[(4'hb):(4'h8)]) && ((^($signed(reg238) ?
          wire233 : (^wire233))) && reg240));
      reg242 <= $signed(wire233[(1'h1):(1'h1)]);
    end
  always
    @(posedge clk) begin
      reg243 <= (($signed((!(wire236 ? wire235 : reg239))) ?
              (($unsigned(reg242) ?
                  (reg239 & wire233) : (wire236 <<< wire234)) || wire235[(4'he):(3'h4)]) : reg241[(2'h2):(1'h0)]) ?
          ((wire236 ?
              wire236 : $signed(wire236)) ^~ (reg238[(3'h5):(2'h3)] << {$signed((8'ha1))})) : (+$signed(($unsigned(reg238) & $unsigned(reg240)))));
      for (forvar244 = (1'h0); (forvar244 < (1'h1)); forvar244 = (forvar244 + (1'h1)))
        begin
          reg245 <= (forvar244[(4'hd):(4'h8)] ?
              $signed(({$unsigned(reg243)} < forvar244[(3'h5):(2'h3)])) : (~&$signed((~^wire237[(3'h4):(1'h0)]))));
          reg246 = ($unsigned(((&(reg238 << reg241)) ?
                  wire237 : $unsigned(reg239[(3'h6):(3'h5)]))) ?
              ((($unsigned(forvar244) <<< (reg242 ?
                      reg243 : (8'haa))) ^~ ($signed(reg238) <<< $signed(reg243))) ?
                  $unsigned(forvar244) : wire233) : $unsigned((+$unsigned($unsigned(reg239)))));
        end
    end
  assign wire247 = reg239[(3'h7):(3'h5)];
  always
    @(posedge clk) begin
      reg248 <= wire235;
      reg249 <= (reg243 ?
          reg248[(2'h3):(2'h3)] : ((~^$unsigned({wire235})) ?
              (reg238[(3'h5):(2'h2)] > $unsigned($unsigned(reg240))) : (^{(-wire247),
                  $unsigned(reg245)})));
      for (forvar250 = (1'h0); (forvar250 < (2'h3)); forvar250 = (forvar250 + (1'h1)))
        begin
          reg251 <= (|(8'h9f));
          for (forvar252 = (1'h0); (forvar252 < (1'h1)); forvar252 = (forvar252 + (1'h1)))
            begin
              reg253 <= $unsigned($unsigned($unsigned((&(+wire236)))));
              reg254 <= (((($signed((8'ha1)) ?
                  (~^forvar244) : {reg251}) & (~^$signed(reg245))) << reg251) <= (~wire247[(3'h6):(2'h2)]));
            end
          reg255 <= $signed($signed((reg246[(4'h8):(1'h0)] ~^ {(reg253 << reg254),
              $signed(reg249)})));
          reg256 <= $signed({reg240});
          reg257 <= ($signed({(forvar250 ?
                  $unsigned(reg241) : (reg255 ~^ reg251))}) <= $unsigned(wire233));
        end
      reg258 = wire237;
    end
  assign wire259 = reg248[(4'h8):(1'h1)];
  always
    @(posedge clk) begin
      reg260 <= $unsigned({$signed(wire236), (~$signed((reg253 <= reg256)))});
      reg261 <= (+$signed(reg243));
    end
  always
    @(posedge clk) begin
      reg262 = {$signed(reg242[(2'h3):(2'h2)]), reg260};
      reg263 = ({wire237[(3'h7):(3'h7)]} && (-reg243[(4'h8):(1'h1)]));
      reg264 = (8'hb3);
      reg265 <= ({(8'ha6), (^~$unsigned({(8'hb0)}))} ?
          reg246 : $unsigned((((+(7'h42)) ? (&reg248) : (^~(8'ha3))) ?
              reg263 : ($signed(reg241) != $signed(reg241)))));
      reg266 <= $unsigned(wire259);
    end
  always
    @(posedge clk) begin
      for (forvar267 = (1'h0); (forvar267 < (2'h2)); forvar267 = (forvar267 + (1'h1)))
        begin
          for (forvar268 = (1'h0); (forvar268 < (1'h0)); forvar268 = (forvar268 + (1'h1)))
            begin
              reg269 <= reg253;
              reg270 <= $signed((~$unsigned((8'hb8))));
              reg271 = reg263[(3'h6):(2'h3)];
              reg272 <= $unsigned(($signed($signed(reg243[(3'h4):(3'h4)])) > $unsigned(((+forvar244) ^~ (8'hbc)))));
            end
          for (forvar273 = (1'h0); (forvar273 < (2'h2)); forvar273 = (forvar273 + (1'h1)))
            begin
              reg274 <= reg254[(2'h3):(1'h0)];
              reg275 <= $signed((~^(reg270 ?
                  ($unsigned(wire237) ?
                      (+reg253) : $unsigned(reg260)) : forvar273)));
              reg276 <= wire233[(3'h7):(3'h4)];
            end
        end
      reg277 <= (~&reg275[(2'h2):(2'h2)]);
      reg278 = wire237;
      reg279 <= $unsigned(wire247);
    end
  always
    @(posedge clk) begin
      reg280 <= $unsigned((~^reg239[(3'h5):(1'h1)]));
      reg281 <= {reg277, (reg256[(3'h4):(3'h4)] ? reg246 : wire235)};
      reg282 <= reg262[(1'h1):(1'h0)];
    end
  always
    @(posedge clk) begin
      for (forvar283 = (1'h0); (forvar283 < (1'h0)); forvar283 = (forvar283 + (1'h1)))
        begin
          reg284 <= (reg282[(2'h2):(1'h0)] ?
              (reg254 ?
                  $signed(reg265[(2'h3):(2'h2)]) : reg246) : ((reg271 > reg279[(3'h5):(3'h4)]) ?
                  reg260 : wire235));
          reg285 <= $unsigned(reg253[(3'h7):(2'h3)]);
          reg286 <= $unsigned((({(reg251 ? reg262 : reg277), {reg274}} ?
              reg256 : $signed((wire234 ?
                  reg270 : reg263))) ~^ $unsigned({$unsigned(reg272),
              {reg265}})));
        end
      reg287 <= (((|$unsigned(((8'hbe) == reg278))) ?
              {(reg245[(4'h9):(4'h9)] ~^ reg254[(3'h4):(2'h2)]),
                  reg258} : reg279[(3'h5):(2'h3)]) ?
          (($signed($signed((8'hbc))) ?
              ($signed(forvar250) <<< reg279[(1'h0):(1'h0)]) : wire237) >= $signed($signed((~wire237)))) : $unsigned((7'h42)));
      reg288 <= wire236[(2'h2):(2'h2)];
      for (forvar289 = (1'h0); (forvar289 < (1'h0)); forvar289 = (forvar289 + (1'h1)))
        begin
          reg290 <= (8'hbb);
          reg291 <= $unsigned(((|(~|(reg284 >> reg245))) ?
              (-(reg242 ? reg279 : $unsigned(reg286))) : (&$signed({reg246}))));
          reg292 = reg260;
          reg293 <= (!$signed(wire236));
          for (forvar294 = (1'h0); (forvar294 < (2'h3)); forvar294 = (forvar294 + (1'h1)))
            begin
              reg295 <= ((wire247 <= (8'hb3)) ?
                  $unsigned($signed(($unsigned(forvar273) | (~|reg258)))) : (7'h44));
              reg296 <= (~^$unsigned(reg266[(5'h10):(4'h9)]));
              reg297 <= (|{reg249, reg257[(2'h3):(2'h2)]});
            end
        end
    end
  assign wire298 = reg255;
  always
    @(posedge clk) begin
      for (forvar299 = (1'h0); (forvar299 < (2'h2)); forvar299 = (forvar299 + (1'h1)))
        begin
          reg300 <= $unsigned((({(+reg246)} > $signed((reg287 != forvar267))) ?
              (+$signed(reg260[(3'h5):(1'h0)])) : reg239[(4'ha):(2'h3)]));
          reg301 <= reg297[(1'h0):(1'h0)];
          reg302 <= forvar268[(3'h5):(2'h2)];
          reg303 <= $signed(reg274[(3'h7):(3'h4)]);
        end
    end
  always
    @(posedge clk) begin
      reg304 <= reg272[(4'hd):(2'h2)];
      reg305 <= wire235;
      reg306 <= reg297[(3'h7):(1'h1)];
      reg307 = ($signed(((reg295[(3'h7):(1'h0)] ? reg255 : $signed((8'hbe))) ?
              (~^$unsigned(reg287)) : ((~|reg264) >> $signed(reg251)))) ?
          wire237 : ({($unsigned(wire234) ?
                  reg253 : $unsigned(wire259))} | $signed({((8'h9f) * reg245),
              $signed((8'ha4))})));
      reg308 = reg286[(4'hb):(4'hb)];
    end
  assign wire309 = (~|$signed(wire235));
  always
    @(posedge clk) begin
      reg310 = $signed($unsigned($unsigned(((~&reg253) ?
          (reg265 ? (8'ha0) : reg302) : $unsigned((8'h9d))))));
      reg311 = ({(reg257 ~^ reg284[(3'h4):(2'h3)])} ?
          $signed($unsigned($signed((reg270 ?
              reg266 : reg285)))) : ((reg307[(1'h1):(1'h1)] <= (8'ha9)) > $unsigned(reg305)));
    end
  assign wire312 = ((~&(reg310[(2'h2):(2'h2)] ?
                           (reg301[(1'h1):(1'h0)] ?
                               $signed(wire236) : forvar252) : ($signed(reg288) + wire298))) ?
                       (!(8'h9f)) : (reg270[(2'h3):(1'h0)] >>> (^~(&(reg293 > reg287)))));
  always
    @(posedge clk) begin
      for (forvar313 = (1'h0); (forvar313 < (2'h3)); forvar313 = (forvar313 + (1'h1)))
        begin
          reg314 = reg278;
          if (reg282)
            begin
              reg315 <= forvar268[(1'h1):(1'h1)];
            end
          else
            begin
              reg315 <= reg285[(4'hc):(4'h9)];
              reg316 <= ((reg311[(2'h2):(1'h0)] ~^ {(reg239[(4'ha):(4'ha)] == (!reg265))}) ?
                  reg270 : (^~$signed($unsigned($signed(forvar294)))));
              reg317 = $unsigned((({reg258[(3'h4):(3'h4)]} ?
                      ({reg239, reg288} ?
                          wire259 : (reg297 ?
                              (8'ha0) : reg256)) : (reg251[(2'h3):(2'h3)] ?
                          $signed(reg281) : $signed(reg315))) ?
                  (~|($signed(reg249) ?
                      (^wire259) : (|reg242))) : {($signed((8'ha2)) ?
                          $signed(forvar250) : $signed(reg238))}));
              reg318 = (reg258[(2'h2):(2'h2)] ?
                  $unsigned(({{reg253}, (reg264 == reg291)} >> {(~^reg301),
                      {reg292,
                          reg290}})) : $unsigned((^((|reg242) << forvar273))));
              reg319 <= $signed({(~&(reg238 ~^ $unsigned(reg256)))});
            end
          reg320 <= (forvar283[(2'h3):(2'h3)] <= $unsigned(reg319));
          for (forvar321 = (1'h0); (forvar321 < (1'h0)); forvar321 = (forvar321 + (1'h1)))
            begin
              reg322 <= $signed((~|($unsigned((reg243 ? reg282 : (7'h41))) ?
                  $unsigned(reg238) : ((reg238 >> reg286) != forvar250))));
            end
          reg323 <= wire312[(1'h0):(1'h0)];
        end
      reg324 <= ((($unsigned($unsigned(reg264)) ?
              $signed($unsigned(reg288)) : {(reg291 & forvar273)}) && {reg319,
              $signed((reg271 || reg318))}) ?
          (reg318[(3'h4):(2'h2)] >> (forvar244 ?
              (~&reg301[(2'h3):(1'h1)]) : $unsigned({wire234,
                  reg307}))) : $signed((8'h9c)));
    end
  always
    @(posedge clk) begin
      for (forvar325 = (1'h0); (forvar325 < (3'h4)); forvar325 = (forvar325 + (1'h1)))
        begin
          reg326 <= (~|((^((-(8'hbe)) ?
                  (reg249 ~^ (8'hba)) : reg255[(2'h3):(2'h3)])) ?
              (~&reg248) : ((~|forvar299) + ((+reg248) ?
                  $signed(forvar313) : $unsigned(reg304)))));
          reg327 <= reg241;
          reg328 <= {(&$signed($unsigned({wire233, reg253}))),
              (+$signed((~^(&reg253))))};
        end
      reg329 <= ((~$unsigned(reg284[(4'h9):(1'h0)])) ?
          reg292[(5'h12):(4'h8)] : $unsigned(reg308[(2'h3):(2'h2)]));
      reg330 = reg301;
      reg331 <= reg277[(1'h1):(1'h0)];
      reg332 <= (7'h42);
    end
  always
    @(posedge clk) begin
      reg333 <= ($unsigned(reg249) * $signed(wire312[(1'h1):(1'h1)]));
      reg334 = (!$signed({$unsigned(wire236)}));
    end
  always
    @(posedge clk) begin
      reg335 <= (reg315[(5'h12):(3'h6)] ? reg285[(4'h9):(1'h0)] : reg286);
      reg336 <= (|reg290);
      reg337 <= {reg270[(2'h3):(2'h3)]};
    end
  always
    @(posedge clk) begin
      reg338 <= ({$signed(reg303)} <<< (~|$unsigned((+reg248[(2'h2):(2'h2)]))));
      reg339 = ((wire312[(1'h0):(1'h0)] ?
              reg337[(2'h2):(1'h0)] : reg330[(2'h3):(1'h0)]) ?
          (8'hb6) : ($signed(reg266) ?
              ((8'h9d) > ((reg305 ? reg336 : reg332) ?
                  ((8'hb1) ?
                      (8'hab) : forvar252) : reg256[(2'h3):(2'h3)])) : $unsigned(($unsigned((8'h9c)) ?
                  forvar252[(1'h0):(1'h0)] : reg269[(1'h1):(1'h0)]))));
      reg340 <= reg241[(2'h2):(1'h0)];
      reg341 <= $unsigned(($unsigned(wire233[(1'h0):(1'h0)]) | $unsigned(reg286[(4'he):(4'h9)])));
      for (forvar342 = (1'h0); (forvar342 < (2'h3)); forvar342 = (forvar342 + (1'h1)))
        begin
          reg343 <= $unsigned((reg296 ?
              $signed(reg291[(4'ha):(3'h6)]) : reg324[(3'h4):(2'h3)]));
          reg344 <= $unsigned($unsigned(reg308[(4'ha):(3'h7)]));
          reg345 <= reg311[(5'h11):(3'h5)];
          reg346 <= $signed({reg293[(1'h0):(1'h0)], (8'hab)});
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module688
#( parameter param752 = ({((((8'ha9) ? (8'h9e) : (7'h42)) ? ((8'hab) >> (8'ha5)) : (^(7'h43))) + (((8'ha3) ? (8'ha8) : (8'hb7)) > (^~(8'hbc))))} > ((+(~((8'hb9) + (8'h9d)))) * ((((8'hbd) ~^ (8'hbe)) < (8'ha4)) ? (8'hb5) : ((|(8'hb8)) && (^(8'ha7))))))
, parameter param753 = (((8'hbf) >>> {(param752 ? (~^param752) : (param752 ? param752 : param752)), ((|(8'hbd)) ^~ (param752 <<< (8'ha1)))}) ? ((((&param752) & {param752}) | (+(^param752))) ? param752 : {param752}) : (|(~|(~(param752 >> (8'ha7)))))) )
(y, clk, wire689, wire690, wire691, wire692, wire693);
  output wire [(32'hb1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hc):(1'h0)] wire689;
  input wire signed [(3'h4):(1'h0)] wire690;
  input wire [(3'h6):(1'h0)] wire691;
  input wire [(5'h14):(1'h0)] wire692;
  input wire signed [(5'h10):(1'h0)] wire693;
  wire [(4'he):(1'h0)] wire694;
  wire signed [(3'h4):(1'h0)] wire695;
  reg signed [(3'h6):(1'h0)] reg696 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg697 = (1'h0);
  reg [(4'hc):(1'h0)] reg698 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire699;
  reg [(4'hb):(1'h0)] forvar700 = (1'h0);
  reg [(4'h8):(1'h0)] reg701 = (1'h0);
  reg [(4'h8):(1'h0)] reg702 = (1'h0);
  reg [(4'hd):(1'h0)] reg703 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg704 = (1'h0);
  reg [(4'he):(1'h0)] reg705 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire706;
  reg signed [(3'h7):(1'h0)] reg707 = (1'h0);
  wire signed [(4'he):(1'h0)] wire750;
  assign y = {wire694,
                 wire695,
                 reg696,
                 reg697,
                 reg698,
                 wire699,
                 forvar700,
                 reg701,
                 reg702,
                 reg703,
                 reg704,
                 reg705,
                 wire706,
                 reg707,
                 wire750,
                 (1'h0)};
  assign wire694 = (($unsigned(wire690[(2'h3):(2'h2)]) ?
                           $signed(wire692) : $unsigned(wire691)) ?
                       ((($signed(wire692) <<< (wire692 <= wire692)) ?
                           wire689 : $unsigned({wire693})) || (wire693 ?
                           $unsigned((wire692 > wire693)) : ((~wire690) ?
                               wire690[(1'h0):(1'h0)] : (~&wire693)))) : wire692[(3'h5):(3'h4)]);
  assign wire695 = ((|wire693) ^~ wire691);
  always
    @(posedge clk) begin
      reg696 <= $signed((($signed($signed(wire692)) ?
              $signed(wire694) : ({wire693, wire692} > wire694)) ?
          wire689 : $signed(wire695[(1'h0):(1'h0)])));
      reg697 <= reg696[(3'h6):(3'h4)];
      reg698 <= $signed(((wire689[(2'h2):(1'h1)] || wire690[(2'h3):(2'h3)]) ?
          {$unsigned($unsigned((8'hbb)))} : ({wire692} ?
              $signed({reg697, wire693}) : $signed($signed((8'ha0))))));
    end
  assign wire699 = (((-wire691[(3'h6):(3'h4)]) != ($unsigned($signed(wire691)) ?
                           $unsigned((wire695 ?
                               wire689 : reg697)) : $signed({wire692,
                               reg697}))) ?
                       $unsigned($unsigned(reg698)) : reg697);
  always
    @(posedge clk) begin
      for (forvar700 = (1'h0); (forvar700 < (2'h3)); forvar700 = (forvar700 + (1'h1)))
        begin
          reg701 <= wire691[(1'h1):(1'h1)];
          reg702 <= (~$unsigned((&$signed(reg698))));
          reg703 <= (~&(|(({wire689, reg698} >> $signed((8'hb2))) ?
              reg697[(1'h1):(1'h0)] : wire694)));
          reg704 <= {(~$unsigned(reg703)),
              ({reg697[(2'h3):(1'h1)], wire699} ?
                  reg696 : $signed(($unsigned(wire699) < $signed(wire691))))};
          reg705 <= $unsigned($unsigned(($signed({reg698,
              (8'hbe)}) <<< wire691[(1'h0):(1'h0)])));
        end
    end
  assign wire706 = (~reg696);
  always
    @(posedge clk) begin
      reg707 <= wire689[(4'h8):(2'h3)];
    end
  module708 modinst751 (wire750, clk, wire692, forvar700, wire706, reg696, reg697);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module533
#( parameter param648 = (-({(((7'h43) != (8'hb2)) ? (8'haa) : ((8'haf) != (8'hb9)))} || (-((7'h44) ? (~^(8'hbf)) : ((8'hb3) ? (8'hb2) : (7'h43)))))) )
(y, clk, wire534, wire535, wire536, wire537, wire538);
  output wire [(32'h203):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire534;
  input wire signed [(5'h15):(1'h0)] wire535;
  input wire [(5'h15):(1'h0)] wire536;
  input wire signed [(4'hd):(1'h0)] wire537;
  input wire signed [(4'ha):(1'h0)] wire538;
  wire signed [(5'h14):(1'h0)] wire647;
  reg signed [(4'hf):(1'h0)] reg646 = (1'h0);
  reg [(4'hc):(1'h0)] reg539 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar540 = (1'h0);
  reg [(4'hd):(1'h0)] reg541 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg542 = (1'h0);
  reg [(4'h9):(1'h0)] reg543 = (1'h0);
  reg [(3'h5):(1'h0)] reg544 = (1'h0);
  reg [(4'hd):(1'h0)] forvar545 = (1'h0);
  reg [(5'h11):(1'h0)] reg546 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg547 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg548 = (1'h0);
  reg [(4'he):(1'h0)] reg549 = (1'h0);
  reg [(3'h7):(1'h0)] reg550 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg551 = (1'h0);
  reg [(3'h6):(1'h0)] reg552 = (1'h0);
  reg [(4'h9):(1'h0)] reg553 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire554;
  reg signed [(3'h4):(1'h0)] reg555 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg556 = (1'h0);
  reg signed [(4'he):(1'h0)] reg557 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar558 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg559 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg560 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg561 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg562 = (1'h0);
  wire [(5'h15):(1'h0)] wire563;
  reg [(5'h10):(1'h0)] reg564 = (1'h0);
  reg [(5'h15):(1'h0)] reg565 = (1'h0);
  reg [(3'h5):(1'h0)] reg566 = (1'h0);
  reg [(4'hb):(1'h0)] forvar567 = (1'h0);
  reg [(5'h14):(1'h0)] forvar568 = (1'h0);
  reg [(3'h6):(1'h0)] reg569 = (1'h0);
  reg [(5'h10):(1'h0)] reg570 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg571 = (1'h0);
  reg [(3'h6):(1'h0)] reg572 = (1'h0);
  reg [(5'h12):(1'h0)] reg573 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg574 = (1'h0);
  reg [(5'h12):(1'h0)] reg575 = (1'h0);
  reg [(4'h9):(1'h0)] reg576 = (1'h0);
  wire [(5'h12):(1'h0)] wire644;
  assign y = {wire647,
                 reg646,
                 reg539,
                 forvar540,
                 reg541,
                 reg542,
                 reg543,
                 reg544,
                 forvar545,
                 reg546,
                 reg547,
                 reg548,
                 reg549,
                 reg550,
                 reg551,
                 reg552,
                 reg553,
                 wire554,
                 reg555,
                 reg556,
                 reg557,
                 forvar558,
                 reg559,
                 reg560,
                 reg561,
                 reg562,
                 wire563,
                 reg564,
                 reg565,
                 reg566,
                 forvar567,
                 forvar568,
                 reg569,
                 reg570,
                 reg571,
                 reg572,
                 reg573,
                 reg574,
                 reg575,
                 reg576,
                 wire644,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg539 <= ($signed($unsigned(($unsigned(wire534) >> (wire534 << wire537)))) <= wire536[(1'h1):(1'h1)]);
      for (forvar540 = (1'h0); (forvar540 < (2'h2)); forvar540 = (forvar540 + (1'h1)))
        begin
          reg541 <= wire534;
          reg542 <= ((wire538 | (wire536[(5'h15):(5'h15)] >>> wire538)) ?
              $signed(wire538) : $signed($signed(wire536)));
          reg543 = (reg541[(2'h2):(2'h2)] <= (reg539 ? wire534 : reg542));
        end
      reg544 <= {(wire536 >>> $signed(((reg539 >>> reg539) ?
              (wire538 + reg542) : $unsigned(wire537)))),
          ((|((-reg541) ? $unsigned(wire534) : (8'hb6))) ?
              ((^{(8'hac), reg541}) ?
                  $unsigned(forvar540[(2'h2):(1'h0)]) : wire536) : ($signed($unsigned(forvar540)) ?
                  (8'ha4) : (wire534[(3'h6):(1'h0)] ?
                      (!(8'ha1)) : $signed(reg542))))};
      for (forvar545 = (1'h0); (forvar545 < (3'h4)); forvar545 = (forvar545 + (1'h1)))
        begin
          reg546 = (forvar540 << (|(reg542[(3'h5):(2'h2)] << {reg542,
              $signed(wire534)})));
          reg547 = ($unsigned($unsigned((&reg542[(4'h9):(3'h4)]))) ^ $signed($unsigned(wire536)));
          reg548 <= (~forvar545);
          reg549 = (reg542 ? (8'haf) : forvar540[(1'h0):(1'h0)]);
          reg550 <= (^reg541[(2'h3):(1'h0)]);
        end
    end
  always
    @(posedge clk) begin
      reg551 = $signed((((~(^reg550)) ?
          wire537 : $signed((reg549 ? reg544 : reg539))) <= ((wire538 ?
              (wire538 < wire537) : wire538[(3'h4):(2'h2)]) ?
          (+(wire535 << reg547)) : reg539[(4'hc):(1'h0)])));
      reg552 <= $signed($signed((~&{(wire536 ^ forvar540)})));
    end
  always
    @(posedge clk) begin
      reg553 = reg542[(3'h5):(2'h3)];
    end
  assign wire554 = $signed((~|{$unsigned(((8'hb0) ? (7'h42) : forvar545)),
                       (~forvar540[(1'h1):(1'h0)])}));
  always
    @(posedge clk) begin
      reg555 <= {($signed({$unsigned(reg542), $signed(reg543)}) ?
              $signed((wire535[(1'h1):(1'h0)] ?
                  reg553[(3'h6):(1'h1)] : $unsigned(reg547))) : wire535[(3'h6):(3'h6)]),
          $unsigned(wire535[(3'h5):(2'h3)])};
      reg556 <= reg547[(2'h2):(2'h2)];
      reg557 <= $unsigned(reg553);
      for (forvar558 = (1'h0); (forvar558 < (2'h3)); forvar558 = (forvar558 + (1'h1)))
        begin
          reg559 <= (forvar558 ?
              ($signed($unsigned((~^reg544))) ?
                  ($signed((reg541 ? reg551 : reg551)) ?
                      reg543[(1'h1):(1'h1)] : forvar545[(1'h0):(1'h0)]) : forvar558[(3'h7):(1'h1)]) : $signed(((!(&reg544)) ?
                  reg553[(2'h2):(1'h1)] : (!(reg552 <= reg552)))));
          reg560 <= {wire536};
        end
    end
  always
    @(posedge clk) begin
      reg561 = reg555[(3'h4):(1'h1)];
      reg562 <= $signed((forvar540 & reg544[(2'h3):(1'h0)]));
    end
  assign wire563 = (wire554 ?
                       reg557[(4'ha):(4'ha)] : $signed({(-(reg549 + reg551)),
                           reg547}));
  always
    @(posedge clk) begin
      reg564 <= (!{$signed(reg551),
          ((&((8'hb2) << wire535)) ?
              reg543[(3'h4):(1'h0)] : ((reg559 ?
                  forvar558 : reg562) ^~ $signed(wire563)))});
      reg565 <= (((~^reg552) ~^ (|$unsigned($unsigned(forvar545)))) * $unsigned((({reg547,
                  reg539} ?
              (forvar540 << reg564) : {reg541}) ?
          ($unsigned(reg541) * reg550[(3'h7):(3'h4)]) : ((~&wire554) > ((8'hb2) * reg559)))));
      reg566 <= ((wire554 ~^ ((reg549 ? {reg559, wire535} : (~^wire554)) ?
              ($unsigned(reg547) ? (|reg555) : (reg550 > reg544)) : (7'h40))) ?
          {(reg544[(1'h0):(1'h0)] <<< reg559[(3'h6):(3'h6)]),
              $signed({(reg559 == reg551)})} : $unsigned($unsigned(($unsigned((8'h9f)) || (reg551 ~^ reg552)))));
      for (forvar567 = (1'h0); (forvar567 < (3'h4)); forvar567 = (forvar567 + (1'h1)))
        begin
          for (forvar568 = (1'h0); (forvar568 < (2'h2)); forvar568 = (forvar568 + (1'h1)))
            begin
              reg569 <= (reg542 ?
                  ($unsigned((!$unsigned(wire535))) - $signed(((wire537 ?
                          reg542 : wire538) ?
                      (reg566 ? reg544 : forvar540) : (reg566 ?
                          reg561 : wire538)))) : $unsigned($signed($signed($signed(wire535)))));
              reg570 <= (((8'hba) ?
                  $signed(((reg546 ?
                      wire535 : forvar545) || (8'hb0))) : {reg539[(1'h0):(1'h0)]}) == wire538);
              reg571 <= {(reg560[(5'h10):(3'h4)] ?
                      wire563 : $unsigned($signed(((8'hbe) ?
                          wire535 : reg559))))};
              reg572 <= (~^(($unsigned(reg548[(4'h9):(1'h0)]) >>> (~|$unsigned(wire563))) <= reg542));
            end
          reg573 <= (^(7'h42));
          reg574 = reg573[(3'h5):(2'h3)];
          reg575 <= $signed(reg566);
        end
      reg576 <= wire554;
    end
  module577 modinst645 (wire644, clk, reg565, forvar568, wire537, forvar545, wire535);
  always
    @(posedge clk) begin
      reg646 <= ((reg573[(4'hc):(4'ha)] > reg541) | {(-wire535[(3'h7):(1'h0)])});
    end
  assign wire647 = $unsigned(wire563);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module577  (y, clk, wire582, wire581, wire580, wire579, wire578);
  output wire [(32'h263):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire582;
  input wire signed [(5'h14):(1'h0)] wire581;
  input wire signed [(4'hd):(1'h0)] wire580;
  input wire [(4'hd):(1'h0)] wire579;
  input wire signed [(5'h15):(1'h0)] wire578;
  reg signed [(4'h8):(1'h0)] reg643 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg642 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg641 = (1'h0);
  reg [(3'h4):(1'h0)] reg640 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire639;
  reg signed [(2'h3):(1'h0)] reg638 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg637 = (1'h0);
  reg [(4'h8):(1'h0)] reg636 = (1'h0);
  reg [(4'he):(1'h0)] reg635 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire634;
  wire signed [(4'h8):(1'h0)] wire633;
  wire [(5'h12):(1'h0)] wire632;
  wire [(4'h9):(1'h0)] wire631;
  reg [(4'ha):(1'h0)] reg630 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg629 = (1'h0);
  reg [(5'h15):(1'h0)] reg628 = (1'h0);
  reg [(3'h6):(1'h0)] reg627 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg626 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg625 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg624 = (1'h0);
  reg [(5'h11):(1'h0)] reg623 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg622 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire621;
  reg [(5'h13):(1'h0)] reg620 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg619 = (1'h0);
  reg [(2'h3):(1'h0)] reg618 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg617 = (1'h0);
  reg [(4'h9):(1'h0)] reg616 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg615 = (1'h0);
  reg [(3'h5):(1'h0)] reg614 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire613;
  wire signed [(4'h8):(1'h0)] wire612;
  reg signed [(2'h2):(1'h0)] reg611 = (1'h0);
  reg [(4'he):(1'h0)] reg610 = (1'h0);
  reg [(5'h12):(1'h0)] reg609 = (1'h0);
  reg [(2'h3):(1'h0)] forvar608 = (1'h0);
  reg [(4'hc):(1'h0)] reg607 = (1'h0);
  reg [(2'h2):(1'h0)] reg606 = (1'h0);
  reg [(5'h10):(1'h0)] reg605 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg604 = (1'h0);
  reg [(4'hd):(1'h0)] reg603 = (1'h0);
  reg [(5'h10):(1'h0)] reg602 = (1'h0);
  reg [(3'h4):(1'h0)] reg601 = (1'h0);
  reg [(3'h7):(1'h0)] forvar600 = (1'h0);
  reg [(5'h12):(1'h0)] reg599 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg598 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg597 = (1'h0);
  reg [(4'hc):(1'h0)] reg596 = (1'h0);
  reg [(2'h3):(1'h0)] reg595 = (1'h0);
  reg [(2'h3):(1'h0)] forvar594 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg593 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar592 = (1'h0);
  reg [(4'h8):(1'h0)] reg591 = (1'h0);
  reg [(3'h5):(1'h0)] reg590 = (1'h0);
  reg [(4'hc):(1'h0)] reg589 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg588 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg587 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg586 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg585 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg584 = (1'h0);
  wire [(5'h15):(1'h0)] wire583;
  assign y = {reg643,
                 reg642,
                 reg641,
                 reg640,
                 wire639,
                 reg638,
                 reg637,
                 reg636,
                 reg635,
                 wire634,
                 wire633,
                 wire632,
                 wire631,
                 reg630,
                 reg629,
                 reg628,
                 reg627,
                 reg626,
                 reg625,
                 reg624,
                 reg623,
                 reg622,
                 wire621,
                 reg620,
                 reg619,
                 reg618,
                 reg617,
                 reg616,
                 reg615,
                 reg614,
                 wire613,
                 wire612,
                 reg611,
                 reg610,
                 reg609,
                 forvar608,
                 reg607,
                 reg606,
                 reg605,
                 reg604,
                 reg603,
                 reg602,
                 reg601,
                 forvar600,
                 reg599,
                 reg598,
                 reg597,
                 reg596,
                 reg595,
                 forvar594,
                 reg593,
                 forvar592,
                 reg591,
                 reg590,
                 reg589,
                 reg588,
                 reg587,
                 reg586,
                 reg585,
                 reg584,
                 wire583,
                 (1'h0)};
  assign wire583 = ($signed({wire579, $signed($signed(wire578))}) - wire580);
  always
    @(posedge clk) begin
      reg584 <= (!wire581);
      reg585 <= {reg584[(4'hb):(4'h8)]};
      reg586 = ({(($unsigned(reg585) ? (reg585 || reg584) : {(7'h43), reg584}) ?
                  reg584 : reg585),
              ((8'hbb) == (^~((8'hb0) ? reg585 : wire578)))} ?
          $unsigned((^~reg585)) : $signed($unsigned((reg585 ?
              (8'hbf) : (reg585 >= wire581)))));
      reg587 = (^~{(8'hab)});
    end
  always
    @(posedge clk) begin
      reg588 <= {wire581};
      reg589 = (~wire583[(1'h1):(1'h0)]);
    end
  always
    @(posedge clk) begin
      reg590 <= $unsigned(((8'ha7) ?
          ($signed($signed(wire579)) >>> (8'ha3)) : (($signed(wire583) ?
                  (wire578 ? wire583 : (8'hac)) : {reg584}) ?
              {$unsigned(reg584),
                  wire582[(4'hb):(4'h8)]} : (^wire580[(2'h3):(2'h2)]))));
      reg591 <= ($unsigned($signed({reg588[(2'h2):(1'h1)]})) & (-((~|(reg588 ?
          (8'ha7) : wire581)) >>> $signed(((8'ha3) ? wire583 : wire578)))));
      for (forvar592 = (1'h0); (forvar592 < (2'h2)); forvar592 = (forvar592 + (1'h1)))
        begin
          reg593 = reg591[(2'h2):(1'h0)];
          for (forvar594 = (1'h0); (forvar594 < (1'h1)); forvar594 = (forvar594 + (1'h1)))
            begin
              reg595 <= ($signed($unsigned($unsigned(reg591[(2'h2):(1'h0)]))) - $signed($unsigned(reg585)));
              reg596 <= $unsigned(wire578[(4'h9):(3'h6)]);
              reg597 <= forvar592[(3'h4):(2'h2)];
              reg598 = wire580;
            end
          reg599 <= $signed((!((7'h42) ?
              ((~&forvar592) == $unsigned(wire583)) : {$unsigned(reg589)})));
          for (forvar600 = (1'h0); (forvar600 < (1'h1)); forvar600 = (forvar600 + (1'h1)))
            begin
              reg601 <= wire581[(5'h13):(2'h3)];
            end
          reg602 = ((((~(^wire579)) ?
                  (reg586 && {forvar600}) : ($unsigned(wire578) ?
                      $unsigned(forvar600) : reg597)) <= reg586) ?
              reg599[(5'h10):(1'h0)] : (|reg590));
        end
      reg603 <= $signed($signed($unsigned(reg588[(2'h2):(2'h2)])));
    end
  always
    @(posedge clk) begin
      reg604 = reg593;
      reg605 <= (!($signed($unsigned({reg585})) == (~&reg584[(3'h6):(2'h2)])));
      reg606 <= forvar600;
      reg607 = (reg604 + $signed(($unsigned($signed(reg595)) ^~ $signed($unsigned(reg605)))));
      for (forvar608 = (1'h0); (forvar608 < (1'h1)); forvar608 = (forvar608 + (1'h1)))
        begin
          reg609 <= (((wire581 ?
              (^$signed(reg587)) : (|(reg599 <<< forvar594))) > (wire578[(3'h6):(2'h2)] & reg605)) ~^ $unsigned({(reg590 + (forvar594 <= reg605))}));
          reg610 = $signed(wire578);
          reg611 = $unsigned(((reg604 ?
                  (reg588 || reg597[(4'h9):(3'h6)]) : ($signed(forvar608) ?
                      $unsigned((8'h9e)) : reg610[(4'hb):(4'h8)])) ?
              (~((forvar600 ^ reg610) >= (^reg605))) : (~^((reg588 ?
                  reg603 : reg602) != (reg585 ? forvar608 : reg610)))));
        end
    end
  assign wire612 = {$signed($signed(reg595))};
  assign wire613 = reg590;
  always
    @(posedge clk) begin
      reg614 = {$signed(($signed((~^(8'h9d))) ^ reg584[(3'h6):(2'h2)])),
          reg611};
      reg615 = (forvar592 * reg597);
      reg616 <= (8'hba);
      reg617 <= ((reg604 ?
              (+(reg607[(1'h0):(1'h0)] <<< ((8'hbb) ?
                  reg609 : reg607))) : (^{(&wire579), $unsigned(forvar608)})) ?
          $signed(reg584[(2'h3):(2'h3)]) : reg590[(3'h5):(2'h3)]);
    end
  always
    @(posedge clk) begin
      reg618 <= (^reg590);
      reg619 <= $signed((&(($signed(reg605) == $signed(reg615)) ?
          (~(reg609 | forvar600)) : reg606[(1'h1):(1'h1)])));
      reg620 <= (~&{$unsigned(((reg603 && reg610) ?
              (forvar608 ? wire580 : reg603) : reg588[(1'h1):(1'h0)])),
          ({$unsigned((8'hb8)), $unsigned(reg615)} - (reg585 ?
              (~&reg593) : (!reg609)))});
    end
  assign wire621 = $signed(($unsigned(reg610) & $signed({{reg616},
                       reg607[(2'h3):(2'h2)]})));
  always
    @(posedge clk) begin
      reg622 <= $signed($signed((reg614[(3'h4):(3'h4)] >>> (reg614[(3'h5):(2'h3)] | reg609[(3'h6):(3'h6)]))));
      reg623 <= $signed(((^~reg598) ?
          $unsigned({{reg584, wire613}, reg615}) : reg604));
      if ($unsigned(($unsigned($unsigned((reg623 ?
          reg585 : wire613))) <= $signed((wire578 < $signed(reg589))))))
        begin
          reg624 <= reg585[(4'hf):(4'hf)];
          reg625 <= ($unsigned($unsigned((reg586 ?
              reg589[(2'h2):(1'h1)] : reg587[(2'h3):(1'h1)]))) ~^ wire583);
          reg626 <= reg602[(4'ha):(4'h9)];
          reg627 <= forvar592[(3'h6):(2'h3)];
          reg628 = (7'h44);
        end
      else
        begin
          reg624 <= $unsigned((~{$unsigned((wire583 >> (8'ha7))),
              ((^reg593) - (!reg609))}));
        end
      reg629 = (8'ha5);
      reg630 <= (+$unsigned($signed($signed($unsigned(reg585)))));
    end
  assign wire631 = reg590;
  assign wire632 = (8'haa);
  assign wire633 = reg595;
  assign wire634 = reg615;
  always
    @(posedge clk) begin
      reg635 = ((~|$unsigned((-{forvar600}))) ?
          ((8'haf) ?
              (~(~&(wire582 ~^ (8'ha6)))) : reg626[(2'h3):(1'h0)]) : (8'hb8));
      reg636 = (|(-(reg611 || $unsigned(reg610))));
      reg637 = $signed($signed({$unsigned($unsigned(reg584)), reg596}));
      reg638 <= (wire634[(1'h0):(1'h0)] ?
          $signed((reg618[(2'h3):(1'h0)] ^~ $signed((reg636 <= (7'h41))))) : $unsigned($unsigned(((reg585 ?
              reg615 : (7'h41)) ^ (reg607 ? reg589 : (8'hb7))))));
    end
  assign wire639 = (((8'hb3) ?
                           $signed(reg636[(2'h2):(1'h0)]) : $signed(((reg628 - reg614) ?
                               (reg614 < wire579) : $signed(reg618)))) ?
                       wire580 : (reg598 < reg586));
  always
    @(posedge clk) begin
      reg640 <= {($unsigned(((reg606 ? reg605 : reg627) ?
                  (~^reg606) : (wire632 <= (8'hb0)))) ?
              reg615[(2'h2):(1'h0)] : reg607)};
      reg641 = ($unsigned(wire579[(1'h1):(1'h1)]) ~^ reg617[(1'h1):(1'h0)]);
      reg642 <= wire621[(2'h2):(2'h2)];
      reg643 <= reg596[(4'hc):(2'h2)];
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module708  (y, clk, wire713, wire712, wire711, wire710, wire709);
  output wire [(32'h1bc):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire713;
  input wire signed [(4'hb):(1'h0)] wire712;
  input wire [(4'h9):(1'h0)] wire711;
  input wire signed [(3'h4):(1'h0)] wire710;
  input wire signed [(5'h11):(1'h0)] wire709;
  wire [(5'h10):(1'h0)] wire749;
  reg [(4'hd):(1'h0)] reg748 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg747 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar746 = (1'h0);
  wire [(4'he):(1'h0)] wire745;
  wire [(4'h9):(1'h0)] wire744;
  wire [(4'hc):(1'h0)] wire743;
  reg signed [(4'h8):(1'h0)] reg742 = (1'h0);
  reg [(2'h2):(1'h0)] reg741 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg740 = (1'h0);
  reg [(5'h15):(1'h0)] reg739 = (1'h0);
  reg signed [(4'he):(1'h0)] reg738 = (1'h0);
  reg [(2'h3):(1'h0)] reg737 = (1'h0);
  reg [(5'h15):(1'h0)] forvar736 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg735 = (1'h0);
  reg [(3'h7):(1'h0)] reg734 = (1'h0);
  reg [(5'h13):(1'h0)] reg733 = (1'h0);
  reg [(2'h2):(1'h0)] reg732 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg731 = (1'h0);
  reg [(4'hc):(1'h0)] forvar730 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg729 = (1'h0);
  reg [(4'h8):(1'h0)] forvar728 = (1'h0);
  wire signed [(4'he):(1'h0)] wire727;
  wire signed [(5'h14):(1'h0)] wire726;
  wire [(5'h14):(1'h0)] wire725;
  reg signed [(5'h12):(1'h0)] reg724 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg723 = (1'h0);
  reg [(2'h2):(1'h0)] reg722 = (1'h0);
  reg [(5'h13):(1'h0)] reg721 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar720 = (1'h0);
  reg [(4'hf):(1'h0)] reg719 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire718;
  wire signed [(2'h2):(1'h0)] wire717;
  reg signed [(4'ha):(1'h0)] reg716 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg715 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg714 = (1'h0);
  assign y = {wire749,
                 reg748,
                 reg747,
                 forvar746,
                 wire745,
                 wire744,
                 wire743,
                 reg742,
                 reg741,
                 reg740,
                 reg739,
                 reg738,
                 reg737,
                 forvar736,
                 reg735,
                 reg734,
                 reg733,
                 reg732,
                 reg731,
                 forvar730,
                 reg729,
                 forvar728,
                 wire727,
                 wire726,
                 wire725,
                 reg724,
                 reg723,
                 reg722,
                 reg721,
                 forvar720,
                 reg719,
                 wire718,
                 wire717,
                 reg716,
                 reg715,
                 reg714,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg714 <= (wire709 ^~ ((~^(~|{wire709})) ?
          (($unsigned(wire710) + wire712[(1'h0):(1'h0)]) <<< wire712[(2'h2):(1'h0)]) : (^wire711)));
      reg715 = ({(-(^~((8'ha3) ? wire710 : wire711)))} | wire710);
      reg716 <= $signed((wire710[(1'h0):(1'h0)] - {((wire712 ?
              wire710 : reg715) <<< ((8'ha0) ^~ wire712)),
          $unsigned($signed((8'h9c)))}));
    end
  assign wire717 = wire712[(2'h3):(2'h2)];
  assign wire718 = (^(|{$signed($unsigned((8'ha3)))}));
  always
    @(posedge clk) begin
      reg719 <= $signed(wire711[(3'h4):(2'h3)]);
      for (forvar720 = (1'h0); (forvar720 < (1'h0)); forvar720 = (forvar720 + (1'h1)))
        begin
          reg721 <= (+(+$signed($signed({reg715}))));
        end
      reg722 <= $unsigned(wire709);
      reg723 <= ((8'hbe) ? wire710 : (wire711 >>> (~^wire717)));
      reg724 <= {{$unsigned((8'had)), $signed({$signed(reg719)})}};
    end
  assign wire725 = (-wire709[(4'h9):(3'h4)]);
  assign wire726 = $unsigned({wire717[(2'h2):(2'h2)], wire710});
  assign wire727 = (reg721[(3'h6):(3'h5)] ? reg722 : (&wire717));
  always
    @(posedge clk) begin
      for (forvar728 = (1'h0); (forvar728 < (2'h2)); forvar728 = (forvar728 + (1'h1)))
        begin
          reg729 <= (wire712[(1'h0):(1'h0)] << reg714[(3'h5):(2'h3)]);
          for (forvar730 = (1'h0); (forvar730 < (3'h4)); forvar730 = (forvar730 + (1'h1)))
            begin
              reg731 <= (forvar730[(3'h6):(3'h4)] <<< reg721);
              reg732 = wire713;
              reg733 <= (~^((forvar728[(3'h5):(2'h2)] || (+((8'h9d) >>> reg721))) | $signed($signed(wire712))));
              reg734 <= {{($signed((!forvar720)) + (~^(~^reg716)))}};
              reg735 = wire709;
            end
          for (forvar736 = (1'h0); (forvar736 < (1'h1)); forvar736 = (forvar736 + (1'h1)))
            begin
              reg737 <= wire717[(1'h0):(1'h0)];
              reg738 = $signed($unsigned(($signed(reg724) ?
                  {(^~reg733)} : (!(reg731 ? reg715 : forvar736)))));
              reg739 <= {(&$unsigned(forvar736)), $signed(wire710)};
              reg740 = (~wire726);
            end
        end
      reg741 <= (($signed($signed(reg716[(3'h7):(1'h1)])) ?
              wire712[(3'h6):(3'h6)] : reg731) ?
          forvar730[(3'h7):(2'h3)] : (!reg735[(3'h5):(2'h3)]));
      reg742 <= (^~reg723[(4'hc):(1'h1)]);
    end
  assign wire743 = (((~&$unsigned(wire709)) != $signed($unsigned($unsigned((8'hbe))))) - reg723);
  assign wire744 = ((^reg715) & ($signed(reg735) ?
                       (+(8'ha2)) : {((reg723 ? (8'h9c) : reg734) ?
                               $signed((8'hbc)) : (wire717 > reg737))}));
  assign wire745 = reg735;
  always
    @(posedge clk) begin
      for (forvar746 = (1'h0); (forvar746 < (1'h0)); forvar746 = (forvar746 + (1'h1)))
        begin
          reg747 <= ((^~($unsigned(reg719[(4'hc):(3'h7)]) > reg733[(3'h6):(1'h0)])) ?
              {reg739,
                  $unsigned({$signed(reg715)})} : (!((wire727 != reg721[(5'h11):(4'hb)]) ?
                  (+(reg731 ?
                      reg723 : reg722)) : (+forvar720[(2'h3):(2'h3)]))));
        end
      reg748 <= ({($unsigned({reg719}) ^ (~&(reg735 >= (8'ha5)))),
          (wire717[(1'h1):(1'h0)] <= (wire718 == $signed(reg740)))} ^ (~|{(!(wire744 ?
              wire726 : (8'hbc)))}));
    end
  assign wire749 = ((~&(($unsigned(wire711) * $unsigned(wire743)) ?
                       wire744[(4'h8):(1'h1)] : (8'hbc))) >= ((&$unsigned((reg734 ?
                       reg729 : (8'ha8)))) << ($signed($unsigned(wire717)) - reg729[(5'h13):(4'h8)])));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module846  (y, clk, wire847, wire848, wire849, wire850);
  output wire [(32'h1e3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire847;
  input wire signed [(5'h13):(1'h0)] wire848;
  input wire signed [(5'h13):(1'h0)] wire849;
  input wire [(2'h2):(1'h0)] wire850;
  wire [(4'ha):(1'h0)] wire1376;
  reg signed [(4'hc):(1'h0)] reg851 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg852 = (1'h0);
  reg [(4'hb):(1'h0)] reg853 = (1'h0);
  reg [(5'h15):(1'h0)] reg854 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg855 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg856 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg857 = (1'h0);
  reg [(3'h6):(1'h0)] reg858 = (1'h0);
  reg [(4'hb):(1'h0)] reg859 = (1'h0);
  reg [(4'hd):(1'h0)] forvar860 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg861 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg862 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar863 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg864 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg865 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg866 = (1'h0);
  reg [(5'h13):(1'h0)] reg867 = (1'h0);
  reg [(5'h10):(1'h0)] reg860 = (1'h0);
  wire [(5'h14):(1'h0)] wire1163;
  reg signed [(4'ha):(1'h0)] reg1165 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire1166;
  reg [(5'h15):(1'h0)] reg1167 = (1'h0);
  wire [(3'h4):(1'h0)] wire1316;
  wire signed [(5'h15):(1'h0)] wire1318;
  reg signed [(5'h12):(1'h0)] reg1319 = (1'h0);
  reg [(3'h4):(1'h0)] reg1320 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1321 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1322 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1323 = (1'h0);
  reg [(3'h5):(1'h0)] reg1324 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1325 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1326 = (1'h0);
  wire [(5'h15):(1'h0)] wire1327;
  wire signed [(5'h14):(1'h0)] wire1328;
  wire signed [(4'hf):(1'h0)] wire1374;
  assign y = {wire1376,
                 reg851,
                 reg852,
                 reg853,
                 reg854,
                 reg855,
                 reg856,
                 reg857,
                 reg858,
                 reg859,
                 forvar860,
                 reg861,
                 reg862,
                 forvar863,
                 reg864,
                 reg865,
                 reg866,
                 reg867,
                 reg860,
                 wire1163,
                 reg1165,
                 wire1166,
                 reg1167,
                 wire1316,
                 wire1318,
                 reg1319,
                 reg1320,
                 forvar1321,
                 reg1322,
                 reg1323,
                 reg1324,
                 reg1325,
                 reg1326,
                 wire1327,
                 wire1328,
                 wire1374,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg851 <= wire847[(2'h3):(1'h1)];
      if ($signed(reg851))
        begin
          reg852 <= wire849[(4'hd):(2'h3)];
          reg853 <= reg851;
          reg854 = wire850;
          reg855 <= wire848[(2'h3):(1'h0)];
          reg856 <= $signed((reg851 ?
              reg855[(1'h0):(1'h0)] : reg852[(1'h1):(1'h1)]));
        end
      else
        begin
          reg852 <= reg854[(4'h9):(1'h0)];
          reg853 = wire849[(5'h11):(3'h4)];
          reg854 = ($unsigned($unsigned($unsigned($signed(wire849)))) ?
              $signed({wire848[(3'h4):(2'h2)],
                  ($signed(wire848) * $unsigned(reg852))}) : reg854[(1'h1):(1'h1)]);
          reg855 <= $unsigned(wire849[(3'h7):(1'h0)]);
        end
      reg857 = $signed(reg853);
      reg858 <= ($signed((((^~wire850) ? $signed(wire848) : (~|wire850)) ?
              reg857 : ({wire849, reg854} + $unsigned((8'ha7))))) ?
          (|((wire850[(1'h0):(1'h0)] ?
              $signed((8'hae)) : (8'h9f)) >>> reg851)) : ($signed($signed((reg852 ?
                  reg851 : (8'ha4)))) ?
              $signed($signed(wire849)) : reg852[(2'h3):(1'h1)]));
    end
  always
    @(posedge clk) begin
      reg859 <= ($unsigned(reg853) & ($signed((8'h9f)) <= {((wire849 ?
              reg852 : wire848) * $signed((8'haf)))}));
      if ((^~reg852))
        begin
          for (forvar860 = (1'h0); (forvar860 < (1'h1)); forvar860 = (forvar860 + (1'h1)))
            begin
              reg861 <= {reg857, reg856[(4'ha):(4'h8)]};
              reg862 = reg854;
            end
          for (forvar863 = (1'h0); (forvar863 < (2'h2)); forvar863 = (forvar863 + (1'h1)))
            begin
              reg864 <= (+(^$unsigned(reg856[(5'h14):(4'hb)])));
              reg865 <= $signed(forvar863);
              reg866 = {$signed($unsigned(((reg856 ? forvar863 : (8'had)) ?
                      (forvar863 ? reg854 : wire848) : reg865[(1'h1):(1'h1)]))),
                  ($signed($signed(reg861)) ~^ reg864[(2'h2):(2'h2)])};
              reg867 = $signed(forvar860[(4'h9):(1'h0)]);
            end
        end
      else
        begin
          reg860 <= {$unsigned(forvar863[(1'h0):(1'h0)])};
          reg861 <= $unsigned((~^(((-(8'hac)) >= forvar863) != $signed(wire848[(4'hd):(2'h3)]))));
        end
    end
  module868 modinst1164 (.wire869(wire849), .wire870(reg860), .y(wire1163), .clk(clk), .wire872(reg853), .wire871(wire848));
  always
    @(posedge clk) begin
      reg1165 <= (~|($unsigned((~|$signed(wire847))) ?
          $signed((reg857[(4'ha):(3'h7)] < $signed(forvar860))) : (-$unsigned(reg861))));
    end
  assign wire1166 = (8'hb0);
  always
    @(posedge clk) begin
      reg1167 <= $unsigned(wire848[(5'h12):(3'h6)]);
    end
  module1168 modinst1317 (.wire1172(reg867), .wire1171(reg1165), .wire1170(wire848), .y(wire1316), .clk(clk), .wire1169(reg851));
  assign wire1318 = $unsigned($unsigned(reg854[(3'h4):(1'h0)]));
  always
    @(posedge clk) begin
      reg1319 <= (!reg1167[(3'h5):(1'h1)]);
      reg1320 <= ($signed((((|(8'hbd)) ?
              (reg855 ? reg858 : reg859) : $signed(reg1165)) ^~ (8'h9c))) ?
          (reg859[(1'h0):(1'h0)] ~^ ($signed(wire1163[(5'h12):(5'h10)]) ?
              (reg861[(3'h5):(1'h0)] == (reg1165 ^ (7'h41))) : $unsigned($signed(reg1319)))) : reg861);
      for (forvar1321 = (1'h0); (forvar1321 < (1'h1)); forvar1321 = (forvar1321 + (1'h1)))
        begin
          reg1322 <= $signed(((~wire847[(1'h1):(1'h1)]) ?
              wire850 : (~|(+reg860[(3'h6):(2'h3)]))));
          reg1323 <= (|((wire847[(4'hb):(2'h2)] ?
              $unsigned($signed(reg861)) : $unsigned((reg1320 ?
                  reg861 : forvar863))) <= ((~&(reg1165 ^~ wire848)) ?
              (|$signed(reg866)) : $unsigned((reg851 ? (8'had) : reg1165)))));
          reg1324 <= $signed($signed(((^~reg862) || ((+wire1316) ^ reg862[(2'h2):(2'h2)]))));
        end
      reg1325 <= (reg856 ? forvar860[(1'h0):(1'h0)] : (&$unsigned((8'hb7))));
      reg1326 <= reg851;
    end
  assign wire1327 = $unsigned($signed(((reg1322 ?
                        reg867[(2'h2):(1'h0)] : (wire1316 || wire848)) || $signed((8'hac)))));
  assign wire1328 = ((reg856 ?
                            reg866 : $signed(($signed(reg867) > ((8'hb2) ?
                                (8'h9c) : reg1165)))) ?
                        {wire1316} : ($unsigned($unsigned(reg859[(4'h8):(3'h5)])) & (((~reg860) << (!reg856)) >>> (wire847 >> wire1316[(2'h3):(2'h2)]))));
  module1329 modinst1375 (wire1374, clk, reg865, reg1325, reg856, reg862, reg1319);
  assign wire1376 = (($unsigned((~^wire1327)) ^~ {$unsigned(reg852)}) <= reg855[(4'ha):(2'h3)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1329  (y, clk, wire1334, wire1333, wire1332, wire1331, wire1330);
  output wire [(32'h1bb):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hf):(1'h0)] wire1334;
  input wire [(2'h3):(1'h0)] wire1333;
  input wire [(4'hf):(1'h0)] wire1332;
  input wire [(5'h12):(1'h0)] wire1331;
  input wire [(4'hd):(1'h0)] wire1330;
  wire signed [(3'h6):(1'h0)] wire1373;
  reg signed [(5'h12):(1'h0)] reg1372 = (1'h0);
  reg [(3'h4):(1'h0)] reg1371 = (1'h0);
  reg [(4'he):(1'h0)] reg1370 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1369 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1368 = (1'h0);
  reg [(4'h8):(1'h0)] reg1367 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1366 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1365 = (1'h0);
  reg [(3'h5):(1'h0)] reg1364 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1363 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1362 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1361 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1360 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1359 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1358 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1357 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1356 = (1'h0);
  reg [(5'h13):(1'h0)] reg1355 = (1'h0);
  reg [(2'h2):(1'h0)] reg1354 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1353 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1352 = (1'h0);
  wire [(3'h6):(1'h0)] wire1351;
  wire [(5'h13):(1'h0)] wire1350;
  wire signed [(4'hb):(1'h0)] wire1349;
  wire [(3'h7):(1'h0)] wire1348;
  reg [(4'hf):(1'h0)] reg1347 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1346 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1345 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1344 = (1'h0);
  reg [(3'h6):(1'h0)] reg1343 = (1'h0);
  wire [(4'h9):(1'h0)] wire1342;
  reg signed [(5'h14):(1'h0)] reg1341 = (1'h0);
  reg [(2'h2):(1'h0)] reg1340 = (1'h0);
  reg [(5'h15):(1'h0)] reg1339 = (1'h0);
  wire [(4'ha):(1'h0)] wire1338;
  wire signed [(4'hb):(1'h0)] wire1337;
  reg [(2'h2):(1'h0)] reg1336 = (1'h0);
  reg [(4'he):(1'h0)] reg1335 = (1'h0);
  assign y = {wire1373,
                 reg1372,
                 reg1371,
                 reg1370,
                 reg1369,
                 reg1368,
                 reg1367,
                 forvar1366,
                 reg1365,
                 reg1364,
                 reg1363,
                 reg1362,
                 reg1361,
                 forvar1360,
                 forvar1359,
                 reg1358,
                 reg1357,
                 reg1356,
                 reg1355,
                 reg1354,
                 forvar1353,
                 reg1352,
                 wire1351,
                 wire1350,
                 wire1349,
                 wire1348,
                 reg1347,
                 reg1346,
                 reg1345,
                 reg1344,
                 reg1343,
                 wire1342,
                 reg1341,
                 reg1340,
                 reg1339,
                 wire1338,
                 wire1337,
                 reg1336,
                 reg1335,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1335 <= wire1334;
      reg1336 <= (-wire1332);
    end
  assign wire1337 = $signed((!$signed($unsigned((wire1334 ?
                        wire1332 : wire1332)))));
  assign wire1338 = ((wire1333[(2'h3):(2'h2)] ^ $signed(reg1336)) >> (~((!$unsigned(wire1332)) | ((^wire1333) ?
                        wire1330 : (!reg1336)))));
  always
    @(posedge clk) begin
      reg1339 = (-$unsigned($signed(wire1332[(2'h2):(1'h0)])));
    end
  always
    @(posedge clk) begin
      reg1340 <= reg1336[(1'h0):(1'h0)];
      reg1341 <= $unsigned($unsigned(wire1333));
    end
  assign wire1342 = reg1339;
  always
    @(posedge clk) begin
      reg1343 <= ($unsigned(wire1338) ?
          $signed((7'h44)) : $signed($unsigned((reg1341[(4'hc):(2'h3)] < (reg1336 ?
              wire1337 : (8'hb3))))));
      reg1344 = {({wire1337} << wire1337), $signed((~^$unsigned((~reg1343))))};
      reg1345 <= (reg1341 & $signed(wire1342));
      reg1346 = $signed((~|$signed(($unsigned((8'ha1)) ? (8'ha6) : (8'hb8)))));
      reg1347 <= {(reg1346 != (-(!reg1343[(1'h0):(1'h0)]))), wire1334};
    end
  assign wire1348 = ((((reg1343 ?
                                (&wire1338) : (reg1345 ?
                                    reg1339 : wire1332)) <<< reg1336[(2'h2):(1'h1)]) ?
                            ((|$signed(wire1331)) >>> ((+(8'ha9)) >= $unsigned(wire1332))) : (-$unsigned($unsigned(reg1340)))) ?
                        $signed(($signed((wire1338 ? (8'ha3) : reg1335)) ?
                            $signed($unsigned(wire1330)) : reg1344[(4'h8):(3'h4)])) : reg1339);
  assign wire1349 = ({reg1336[(1'h0):(1'h0)],
                            ($unsigned($unsigned(reg1341)) && {wire1337[(2'h3):(2'h3)],
                                $signed(reg1336)})} ?
                        (+(~&wire1330[(1'h1):(1'h1)])) : (wire1348[(1'h0):(1'h0)] ^~ ($unsigned((reg1343 * (8'hb0))) ^~ $unsigned((wire1334 <<< (8'hbd))))));
  assign wire1350 = ((((reg1341 ? $signed(reg1345) : (&wire1338)) ?
                        $signed((^wire1338)) : reg1346) | (~|(8'ha2))) ~^ reg1344[(3'h6):(3'h5)]);
  assign wire1351 = (&$signed(reg1344));
  always
    @(posedge clk) begin
      reg1352 <= $signed($signed($signed(reg1347)));
      for (forvar1353 = (1'h0); (forvar1353 < (1'h1)); forvar1353 = (forvar1353 + (1'h1)))
        begin
          reg1354 <= (((8'ha4) <= (8'h9e)) ?
              wire1333 : {($unsigned((-reg1340)) <<< {(reg1346 > wire1351),
                      wire1333[(1'h0):(1'h0)]})});
        end
    end
  always
    @(posedge clk) begin
      reg1355 <= {$unsigned((reg1339[(2'h3):(2'h3)] ?
              $unsigned((^~reg1343)) : ({wire1332, reg1344} ?
                  $unsigned(wire1331) : $signed(reg1354)))),
          $signed(((|$unsigned(wire1350)) ^~ wire1338[(3'h5):(2'h3)]))};
      reg1356 <= wire1333;
      reg1357 <= (8'ha3);
      reg1358 <= (((((reg1357 ?
                  reg1347 : (8'ha5)) | $signed(reg1355)) || wire1348) ?
              ({wire1350} ^ (|wire1342)) : $signed($signed(reg1352[(2'h2):(1'h1)]))) ?
          reg1352 : $unsigned($signed((~^(+forvar1353)))));
    end
  always
    @(posedge clk) begin
      for (forvar1359 = (1'h0); (forvar1359 < (2'h3)); forvar1359 = (forvar1359 + (1'h1)))
        begin
          for (forvar1360 = (1'h0); (forvar1360 < (2'h2)); forvar1360 = (forvar1360 + (1'h1)))
            begin
              reg1361 <= ((wire1334 || $signed(((~reg1346) ?
                      (~^wire1332) : (reg1352 < wire1338)))) ?
                  ($unsigned(wire1330[(4'hc):(1'h1)]) <<< (reg1336[(2'h2):(1'h0)] >= ((~^reg1335) | $unsigned(reg1335)))) : wire1333);
              reg1362 <= reg1355;
            end
          reg1363 <= $unsigned((^wire1351[(2'h3):(1'h0)]));
          reg1364 = (&reg1358);
          reg1365 <= $signed($unsigned($signed($signed($unsigned(reg1357)))));
        end
      for (forvar1366 = (1'h0); (forvar1366 < (1'h0)); forvar1366 = (forvar1366 + (1'h1)))
        begin
          reg1367 <= reg1364;
          reg1368 <= ((({(reg1361 < wire1333)} * ($unsigned(wire1349) ^ $signed(reg1365))) >> (8'hbc)) ?
              $signed((~|(8'hb4))) : $signed(($signed((reg1335 & wire1338)) ?
                  $unsigned((wire1330 ? wire1350 : wire1342)) : {(wire1331 ?
                          reg1336 : reg1358),
                      $unsigned((8'hbe))})));
          reg1369 <= (!(8'h9c));
        end
      reg1370 <= ($signed((~|reg1340[(1'h1):(1'h0)])) - reg1340);
      reg1371 <= $signed({$signed((reg1367 ? (~reg1364) : $signed(reg1363))),
          wire1337[(2'h3):(2'h2)]});
    end
  always
    @(posedge clk) begin
      reg1372 <= (wire1351 ^~ wire1332[(1'h1):(1'h0)]);
    end
  assign wire1373 = wire1351;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1168
#( parameter param1315 = ({(-(((7'h43) || (8'hb2)) || (8'hb0))), ((((8'ha6) > (8'hac)) ? ((8'hbb) + (8'had)) : ((8'hac) ? (8'h9f) : (8'ha4))) ? ((8'ha9) ^ {(8'hb0)}) : (((8'hb3) == (8'hbc)) + ((8'haf) && (8'ha3))))} ~^ {((-{(7'h42)}) ? (8'hbd) : (((8'haf) ? (8'ha0) : (8'hb4)) * ((8'hb3) != (8'ha2))))}) )
(y, clk, wire1169, wire1170, wire1171, wire1172);
  output wire [(32'h15e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h9):(1'h0)] wire1169;
  input wire [(3'h4):(1'h0)] wire1170;
  input wire [(2'h3):(1'h0)] wire1171;
  input wire [(5'h13):(1'h0)] wire1172;
  reg [(5'h11):(1'h0)] reg1314 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1313 = (1'h0);
  reg [(4'h8):(1'h0)] reg1312 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1311 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1310 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1309 = (1'h0);
  wire [(3'h4):(1'h0)] wire1308;
  reg [(3'h7):(1'h0)] reg1307 = (1'h0);
  wire [(3'h7):(1'h0)] wire1306;
  reg signed [(4'h9):(1'h0)] reg1305 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1304 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire1302;
  reg signed [(4'h9):(1'h0)] reg1247 = (1'h0);
  reg [(4'hc):(1'h0)] reg1246 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1245 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1244 = (1'h0);
  wire [(3'h7):(1'h0)] wire1243;
  reg [(4'ha):(1'h0)] reg1173 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1174 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1175 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1176 = (1'h0);
  reg [(4'hc):(1'h0)] reg1177 = (1'h0);
  reg [(4'he):(1'h0)] reg1178 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1179 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1180 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1181 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1182 = (1'h0);
  reg [(5'h14):(1'h0)] reg1183 = (1'h0);
  reg [(4'he):(1'h0)] reg1184 = (1'h0);
  wire [(3'h7):(1'h0)] wire1185;
  wire signed [(4'h9):(1'h0)] wire1241;
  assign y = {reg1314,
                 reg1313,
                 reg1312,
                 reg1311,
                 forvar1310,
                 reg1309,
                 wire1308,
                 reg1307,
                 wire1306,
                 reg1305,
                 reg1304,
                 wire1302,
                 reg1247,
                 reg1246,
                 reg1245,
                 forvar1244,
                 wire1243,
                 reg1173,
                 forvar1174,
                 forvar1175,
                 reg1176,
                 reg1177,
                 reg1178,
                 reg1179,
                 reg1180,
                 reg1181,
                 reg1182,
                 reg1183,
                 reg1184,
                 wire1185,
                 wire1241,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1173 <= wire1170;
      for (forvar1174 = (1'h0); (forvar1174 < (1'h1)); forvar1174 = (forvar1174 + (1'h1)))
        begin
          for (forvar1175 = (1'h0); (forvar1175 < (2'h3)); forvar1175 = (forvar1175 + (1'h1)))
            begin
              reg1176 <= (-(~|($signed(forvar1174[(3'h5):(1'h0)]) ?
                  (wire1169 >> $unsigned(forvar1175)) : ($signed(wire1171) & (~^wire1170)))));
              reg1177 <= $signed(forvar1175);
              reg1178 <= (8'ha3);
            end
          reg1179 <= $unsigned({$unsigned(reg1177[(1'h0):(1'h0)]),
              $signed(reg1177)});
        end
    end
  always
    @(posedge clk) begin
      reg1180 <= forvar1175;
      reg1181 <= wire1172[(4'hd):(4'ha)];
      reg1182 <= {$signed(reg1180)};
      reg1183 <= $unsigned((+{(reg1177 >> $signed(reg1178)),
          $unsigned($signed(wire1172))}));
      reg1184 <= {$unsigned(($signed((~forvar1174)) ?
              ((wire1169 ? reg1179 : reg1179) ?
                  (reg1183 + wire1171) : wire1169) : (~^$unsigned(reg1173)))),
          $signed({((~(8'hae)) ?
                  $unsigned(reg1179) : reg1178[(4'h8):(2'h3)])})};
    end
  assign wire1185 = wire1170[(1'h0):(1'h0)];
  module1186 modinst1242 (.wire1190(reg1180), .y(wire1241), .wire1189(reg1182), .wire1191(wire1172), .wire1187(wire1170), .clk(clk), .wire1188(reg1179));
  assign wire1243 = $unsigned(reg1178[(2'h3):(1'h1)]);
  always
    @(posedge clk) begin
      for (forvar1244 = (1'h0); (forvar1244 < (2'h3)); forvar1244 = (forvar1244 + (1'h1)))
        begin
          reg1245 <= (~|(wire1185 ?
              (((~&wire1170) && (^reg1173)) ?
                  (~&(~|forvar1244)) : $unsigned($signed(wire1170))) : $signed((~|(wire1185 ?
                  wire1241 : (8'ha0))))));
          reg1246 <= (^~reg1173);
          reg1247 <= ($unsigned($unsigned($unsigned($unsigned(reg1180)))) >>> ($signed({wire1170[(2'h3):(1'h1)]}) ?
              {((^(8'hae)) ^~ $unsigned(wire1241))} : {(~&(reg1173 ?
                      forvar1244 : forvar1244))}));
        end
    end
  module1248 modinst1303 (.y(wire1302), .wire1249(reg1178), .clk(clk), .wire1251(reg1181), .wire1250(reg1183), .wire1252(forvar1175));
  always
    @(posedge clk) begin
      reg1304 <= $signed(reg1177[(4'hc):(1'h0)]);
      reg1305 <= {wire1169,
          (wire1302 >>> (reg1180 ^~ ((wire1241 ? wire1243 : wire1172) ?
              $unsigned(forvar1174) : $unsigned(wire1172))))};
    end
  assign wire1306 = forvar1174[(2'h2):(1'h1)];
  always
    @(posedge clk) begin
      reg1307 <= $signed((8'h9d));
    end
  assign wire1308 = (reg1177 ?
                        (((|{reg1173, reg1184}) ?
                            wire1169[(4'h8):(4'h8)] : (+wire1243[(3'h4):(2'h2)])) >= ({wire1306[(1'h0):(1'h0)]} ?
                            ((|(8'hb2)) ?
                                $signed(wire1171) : reg1176[(1'h0):(1'h0)]) : ($signed(reg1305) && reg1182[(2'h3):(1'h0)]))) : ($unsigned(reg1173[(2'h2):(1'h0)]) ?
                            (&{$signed(reg1307)}) : reg1183));
  always
    @(posedge clk) begin
      reg1309 = reg1307;
      for (forvar1310 = (1'h0); (forvar1310 < (1'h0)); forvar1310 = (forvar1310 + (1'h1)))
        begin
          reg1311 <= $unsigned(((reg1182[(1'h1):(1'h1)] & {$unsigned((8'haa)),
                  $unsigned(wire1243)}) ?
              $unsigned((^~forvar1175[(1'h0):(1'h0)])) : (forvar1174[(1'h1):(1'h0)] ?
                  ({forvar1174} ?
                      $unsigned((8'hac)) : forvar1175) : (~&reg1177[(3'h7):(1'h1)]))));
        end
      reg1312 = reg1184[(3'h5):(1'h1)];
      reg1313 <= {$unsigned($unsigned((reg1312 ?
              (&wire1185) : $unsigned(forvar1174))))};
      reg1314 <= ((8'h9f) ?
          ((^wire1308) == {{((8'ha7) != (8'hb4))}}) : reg1312);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module868
#( parameter param1162 = ((({((8'hba) ? (7'h44) : (8'hb4)), ((8'h9e) >>> (8'ha1))} ? (((8'hb1) ? (8'h9d) : (7'h40)) ? (~|(8'ha8)) : {(8'hba)}) : (~(!(8'ha8)))) * (~^(((8'hab) ? (8'hb2) : (8'hae)) ^ (~(8'ha7))))) ? (({(^(8'hb2))} ~^ (~^((8'hbe) ? (8'hb7) : (8'hb0)))) ? (-(^{(8'ha5)})) : ((~{(8'hac), (7'h43)}) ? {((8'hab) ? (8'hbf) : (8'h9c)), ((8'h9e) ? (8'hac) : (7'h41))} : ((~^(8'ha9)) << ((8'hb6) ^ (8'h9d))))) : (^((((8'hb4) * (8'hb6)) ^ (7'h43)) ? (((8'ha7) || (8'ha9)) ? ((7'h42) == (8'hb9)) : ((8'hb4) ^ (8'had))) : (!{(8'ha3), (8'ha3)})))) )
(y, clk, wire872, wire871, wire870, wire869);
  output wire [(32'h3b2):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hb):(1'h0)] wire872;
  input wire signed [(5'h13):(1'h0)] wire871;
  input wire signed [(5'h10):(1'h0)] wire870;
  input wire [(5'h12):(1'h0)] wire869;
  reg [(3'h7):(1'h0)] reg1161 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1160 = (1'h0);
  reg [(5'h13):(1'h0)] reg1159 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1158 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1157 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1156 = (1'h0);
  reg [(4'h8):(1'h0)] reg1155 = (1'h0);
  reg [(2'h3):(1'h0)] reg1154 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1153 = (1'h0);
  reg [(2'h2):(1'h0)] reg1152 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1151 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1150 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1149 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1148 = (1'h0);
  reg [(5'h15):(1'h0)] reg1147 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1146 = (1'h0);
  reg [(4'ha):(1'h0)] reg1145 = (1'h0);
  reg [(3'h6):(1'h0)] reg1144 = (1'h0);
  reg [(5'h13):(1'h0)] reg1143 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1142 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1141 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1140 = (1'h0);
  reg [(2'h2):(1'h0)] reg1139 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1138 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1137 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1136 = (1'h0);
  reg [(4'h8):(1'h0)] reg1135 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1134 = (1'h0);
  reg [(4'hd):(1'h0)] reg1133 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire1132;
  wire signed [(3'h6):(1'h0)] wire1131;
  reg [(5'h11):(1'h0)] reg1130 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1129 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire1128;
  wire signed [(2'h3):(1'h0)] wire1127;
  reg [(5'h10):(1'h0)] reg1126 = (1'h0);
  reg [(4'hc):(1'h0)] reg1125 = (1'h0);
  reg [(4'hf):(1'h0)] reg1124 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1123 = (1'h0);
  reg [(3'h7):(1'h0)] reg1122 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1121 = (1'h0);
  reg [(4'ha):(1'h0)] reg1120 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1119 = (1'h0);
  reg [(2'h2):(1'h0)] reg1118 = (1'h0);
  reg [(3'h4):(1'h0)] reg1117 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1116 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1115 = (1'h0);
  reg [(2'h2):(1'h0)] reg1114 = (1'h0);
  reg [(5'h13):(1'h0)] reg1113 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1112 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1111 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1110 = (1'h0);
  wire [(5'h11):(1'h0)] wire1108;
  wire [(4'h8):(1'h0)] wire1073;
  reg [(2'h2):(1'h0)] reg1072 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1071 = (1'h0);
  reg [(2'h3):(1'h0)] reg1070 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1069 = (1'h0);
  reg [(4'he):(1'h0)] reg1068 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1067 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1066 = (1'h0);
  reg [(4'ha):(1'h0)] reg1065 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1064 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire935;
  reg signed [(4'hf):(1'h0)] reg880 = (1'h0);
  reg [(5'h10):(1'h0)] reg879 = (1'h0);
  reg signed [(4'he):(1'h0)] reg878 = (1'h0);
  reg [(3'h7):(1'h0)] reg877 = (1'h0);
  reg signed [(4'he):(1'h0)] reg876 = (1'h0);
  reg [(5'h12):(1'h0)] reg875 = (1'h0);
  reg [(5'h12):(1'h0)] forvar874 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar873 = (1'h0);
  wire [(3'h6):(1'h0)] wire982;
  wire [(5'h15):(1'h0)] wire984;
  wire [(2'h3):(1'h0)] wire985;
  reg signed [(4'ha):(1'h0)] reg986 = (1'h0);
  reg [(3'h7):(1'h0)] reg987 = (1'h0);
  reg [(5'h11):(1'h0)] reg988 = (1'h0);
  reg [(5'h13):(1'h0)] forvar989 = (1'h0);
  reg [(4'he):(1'h0)] reg990 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar991 = (1'h0);
  reg [(4'hb):(1'h0)] reg992 = (1'h0);
  reg [(4'hd):(1'h0)] reg993 = (1'h0);
  wire [(5'h14):(1'h0)] wire1062;
  assign y = {reg1161,
                 reg1160,
                 reg1159,
                 reg1158,
                 forvar1157,
                 reg1156,
                 reg1155,
                 reg1154,
                 reg1153,
                 reg1152,
                 reg1151,
                 reg1150,
                 reg1149,
                 reg1148,
                 reg1147,
                 forvar1146,
                 reg1145,
                 reg1144,
                 reg1143,
                 forvar1142,
                 forvar1141,
                 reg1140,
                 reg1139,
                 reg1138,
                 reg1137,
                 reg1136,
                 reg1135,
                 forvar1134,
                 reg1133,
                 wire1132,
                 wire1131,
                 reg1130,
                 reg1129,
                 wire1128,
                 wire1127,
                 reg1126,
                 reg1125,
                 reg1124,
                 reg1123,
                 reg1122,
                 reg1121,
                 reg1120,
                 reg1119,
                 reg1118,
                 reg1117,
                 reg1116,
                 reg1115,
                 reg1114,
                 reg1113,
                 forvar1112,
                 reg1111,
                 reg1110,
                 wire1108,
                 wire1073,
                 reg1072,
                 reg1071,
                 reg1070,
                 reg1069,
                 reg1068,
                 reg1067,
                 reg1066,
                 reg1065,
                 forvar1064,
                 wire935,
                 reg880,
                 reg879,
                 reg878,
                 reg877,
                 reg876,
                 reg875,
                 forvar874,
                 forvar873,
                 wire982,
                 wire984,
                 wire985,
                 reg986,
                 reg987,
                 reg988,
                 forvar989,
                 reg990,
                 forvar991,
                 reg992,
                 reg993,
                 wire1062,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar873 = (1'h0); (forvar873 < (2'h2)); forvar873 = (forvar873 + (1'h1)))
        begin
          for (forvar874 = (1'h0); (forvar874 < (1'h1)); forvar874 = (forvar874 + (1'h1)))
            begin
              reg875 = $signed((^~($signed($signed(wire869)) >>> forvar873)));
              reg876 <= ($unsigned(forvar874) == (~|(wire870[(1'h1):(1'h0)] ?
                  (((8'h9f) >> wire869) == (~^wire869)) : $unsigned(forvar874))));
              reg877 <= forvar874[(1'h1):(1'h0)];
              reg878 = (&$unsigned($unsigned(wire870)));
            end
          reg879 = reg876[(1'h1):(1'h1)];
          reg880 <= $unsigned(reg878[(2'h3):(1'h0)]);
        end
    end
  module881 modinst936 (wire935, clk, reg880, reg876, reg879, wire871, wire872);
  module937 modinst983 (wire982, clk, reg879, reg880, wire871, wire869);
  assign wire984 = wire872[(2'h2):(1'h1)];
  assign wire985 = forvar874[(5'h11):(4'hc)];
  always
    @(posedge clk) begin
      reg986 <= ((8'ha2) ?
          (8'hb0) : $unsigned((^~(~(reg875 ? wire935 : reg877)))));
      reg987 <= (($signed((-(wire984 - reg875))) ?
          (&(reg880 ?
              (forvar873 ? forvar873 : reg876) : (^~wire872))) : (wire869 ?
              (-$signed(forvar873)) : $unsigned((+reg875)))) | $unsigned((reg986 ?
          {$signed(wire985), (~&wire985)} : ((~&forvar873) ?
              reg875[(2'h2):(1'h0)] : $signed((8'ha8))))));
      reg988 <= reg879;
      for (forvar989 = (1'h0); (forvar989 < (2'h3)); forvar989 = (forvar989 + (1'h1)))
        begin
          reg990 = (~$unsigned(wire872));
          for (forvar991 = (1'h0); (forvar991 < (3'h4)); forvar991 = (forvar991 + (1'h1)))
            begin
              reg992 = $unsigned({(~|wire869[(3'h7):(3'h7)]),
                  (((forvar991 ? forvar874 : reg876) == (forvar991 ?
                          wire984 : wire984)) ?
                      (+(wire984 ? reg988 : (8'ha9))) : {{(8'ha7), reg880}})});
              reg993 <= wire869[(5'h12):(4'h8)];
            end
        end
    end
  module994 modinst1063 (wire1062, clk, reg987, wire870, reg875, wire871, wire935);
  always
    @(posedge clk) begin
      if (wire985[(1'h0):(1'h0)])
        begin
          for (forvar1064 = (1'h0); (forvar1064 < (2'h3)); forvar1064 = (forvar1064 + (1'h1)))
            begin
              reg1065 <= ($signed(forvar873[(2'h3):(2'h3)]) ?
                  ($unsigned((((8'ha4) ?
                      wire935 : reg878) | (~|reg992))) | (({wire982} ?
                      $signed((8'hb5)) : $signed(reg875)) << $unsigned(reg878[(4'ha):(4'h8)]))) : (!$unsigned((^(&forvar1064)))));
              reg1066 <= (reg879[(5'h10):(4'hd)] ?
                  reg875[(5'h10):(4'hf)] : (|({(forvar873 && (8'hbc))} >= $unsigned(wire985[(1'h0):(1'h0)]))));
              reg1067 <= (($unsigned({(+forvar873)}) << $unsigned(reg880[(4'he):(3'h4)])) ~^ (|reg877[(2'h2):(1'h0)]));
              reg1068 <= wire935;
              reg1069 = reg987[(2'h2):(2'h2)];
            end
          reg1070 <= ($signed(forvar874) ?
              wire985 : $unsigned($unsigned({$unsigned(reg876)})));
          reg1071 <= (reg1066 ?
              {reg1070,
                  ($unsigned({wire985,
                      reg986}) | reg876)} : $signed({({reg1066} ?
                      $unsigned(reg876) : (reg879 ? wire871 : forvar989))}));
        end
      else
        begin
          for (forvar1064 = (1'h0); (forvar1064 < (2'h3)); forvar1064 = (forvar1064 + (1'h1)))
            begin
              reg1065 <= reg1070;
              reg1066 = wire870;
              reg1067 <= (($signed(forvar989[(4'h8):(3'h4)]) ?
                  $signed(reg990[(4'h9):(1'h1)]) : $unsigned($signed(((8'had) & (8'ha8))))) - $signed(reg879));
              reg1068 = $unsigned((((forvar989[(4'h9):(2'h3)] ?
                      (^(8'ha9)) : $signed((8'hb2))) ?
                  ($signed(forvar874) * (^~reg1070)) : ((reg990 ?
                          reg1068 : (8'hba)) ?
                      $signed(wire869) : (wire935 <<< reg880))) <<< ($signed($unsigned(reg1067)) ?
                  forvar991 : $signed($unsigned(reg992)))));
              reg1069 <= (&(|wire872[(1'h1):(1'h0)]));
            end
          reg1070 <= (^~(reg875 || (^$unsigned(reg990[(4'h8):(4'h8)]))));
        end
      reg1072 <= reg876[(2'h3):(1'h1)];
    end
  assign wire1073 = (~^reg1069[(2'h2):(1'h0)]);
  module1074 modinst1109 (wire1108, clk, wire1062, wire985, reg1070, wire872);
  always
    @(posedge clk) begin
      reg1110 <= $unsigned($unsigned({(~|$signed(wire872))}));
    end
  always
    @(posedge clk) begin
      reg1111 <= $unsigned((reg877 ?
          (!$signed({reg1070, wire872})) : (wire869[(1'h1):(1'h1)] ?
              $unsigned((forvar874 * reg1068)) : ($unsigned(reg1067) >>> $signed(wire1062)))));
      for (forvar1112 = (1'h0); (forvar1112 < (2'h3)); forvar1112 = (forvar1112 + (1'h1)))
        begin
          reg1113 = wire872;
          if ($unsigned(((8'hac) ?
              $signed(((|wire982) ^~ reg1111[(3'h6):(2'h2)])) : $unsigned($signed(reg990[(2'h2):(1'h0)])))))
            begin
              reg1114 <= ($unsigned(reg1066[(2'h3):(2'h3)]) ?
                  $unsigned((($unsigned(reg1110) ?
                      ((8'hb3) >= reg1067) : (^~reg1065)) * (reg1065[(1'h1):(1'h0)] ~^ (wire985 | reg1068)))) : $unsigned($unsigned(reg1066[(1'h0):(1'h0)])));
              reg1115 = $signed((|($unsigned(reg1067[(4'hd):(4'hc)]) * reg877)));
              reg1116 <= $unsigned($signed({(|$unsigned(reg1111))}));
              reg1117 <= $unsigned(forvar989);
              reg1118 = forvar1064[(2'h3):(2'h3)];
            end
          else
            begin
              reg1114 <= (-(~&forvar1064));
              reg1115 <= ((^~{forvar1064[(3'h4):(1'h0)]}) == $unsigned($unsigned($signed(reg1068))));
            end
          reg1119 <= ((~^$signed($signed(reg880))) ? wire985 : reg1114);
          reg1120 <= (~|(((~^$signed(forvar1112)) - $signed(wire984[(4'hf):(2'h3)])) == (reg878[(1'h0):(1'h0)] << reg993)));
        end
      if (wire1062[(4'hc):(4'hb)])
        begin
          reg1121 <= {((~($unsigned((8'hb6)) == reg1118)) ^~ reg1113[(3'h6):(3'h4)])};
          reg1122 <= $signed($unsigned((^reg1121)));
          reg1123 <= reg1065[(3'h6):(2'h2)];
          reg1124 <= reg1072;
          reg1125 <= $unsigned(((wire982[(3'h5):(1'h0)] * (+wire1062)) ?
              (((-reg875) > ((8'ha5) != reg1065)) > $signed((reg1117 >= reg993))) : wire1108[(4'hd):(4'hd)]));
        end
      else
        begin
          reg1121 = (wire1073[(3'h7):(3'h6)] ^~ (-reg880));
          reg1122 = (reg1065[(3'h5):(2'h2)] ?
              (8'haf) : ($signed(($signed(reg1111) * $signed(reg1120))) ?
                  $signed((~|(reg1113 + wire935))) : reg1125));
          reg1123 = (8'hbc);
          reg1124 <= (~^{(|$unsigned({(7'h42), reg1111})),
              (+reg1069[(2'h3):(1'h0)])});
          reg1125 = ({(reg987[(2'h3):(2'h2)] ?
                  reg880[(4'hf):(4'ha)] : (|(-reg987))),
              reg1120[(4'ha):(1'h0)]} && (-$unsigned({(reg993 ?
                  reg990 : reg1121),
              (8'hbe)})));
        end
      reg1126 <= $unsigned($signed(reg1068));
    end
  assign wire1127 = $signed($signed(((!forvar989) && reg875)));
  assign wire1128 = forvar1112;
  always
    @(posedge clk) begin
      reg1129 <= (((|(&(forvar1112 ? reg875 : reg1114))) ?
              {({wire871, reg878} ?
                      (~|reg878) : $signed((8'hb9)))} : wire982[(1'h1):(1'h0)]) ?
          (((-(8'hb7)) < $signed((~|wire1062))) > ($unsigned({wire982,
              reg1110}) >>> $signed((reg1123 ?
              wire872 : reg1125)))) : (($unsigned((+(8'hb3))) ?
                  wire982[(3'h4):(1'h0)] : ($unsigned((8'hb2)) ?
                      (-wire1062) : $signed(wire872))) ?
              {(reg1118 ? ((8'ha2) >= wire1073) : reg1123[(3'h4):(3'h4)]),
                  {reg1116}} : forvar873));
      reg1130 <= ({reg1072[(1'h0):(1'h0)],
          {$signed($unsigned(wire1073))}} == $unsigned(((~{(7'h42)}) ?
          {reg1129} : ((8'ha7) ? wire1108 : (reg1126 ? (8'ha1) : wire1128)))));
    end
  assign wire1131 = (|({($unsigned((8'h9f)) * reg1068[(1'h1):(1'h1)])} <= ($unsigned(reg992) >>> wire872)));
  assign wire1132 = (+$signed((|wire1127[(1'h1):(1'h0)])));
  always
    @(posedge clk) begin
      reg1133 = $unsigned({(~reg1067[(5'h11):(2'h3)])});
      for (forvar1134 = (1'h0); (forvar1134 < (1'h0)); forvar1134 = (forvar1134 + (1'h1)))
        begin
          reg1135 = (-{reg1070, $unsigned(wire872[(3'h6):(1'h1)])});
        end
    end
  always
    @(posedge clk) begin
      if (reg1071)
        begin
          reg1136 <= {(+($unsigned((reg1124 ?
                  (8'ha8) : forvar873)) ^~ ($signed(forvar991) ?
                  $signed(wire1127) : $unsigned(reg1125)))),
              forvar874[(5'h11):(2'h3)]};
          reg1137 = {$signed((-reg1126[(3'h7):(3'h4)])), reg1115};
        end
      else
        begin
          reg1136 <= $unsigned(reg1065[(4'ha):(4'ha)]);
          reg1137 <= reg986;
          reg1138 <= (+{reg1067[(4'he):(4'hd)]});
          reg1139 <= {$signed($unsigned(((reg1129 ? reg1070 : forvar873) ?
                  $signed((8'ha8)) : reg1137[(4'h9):(1'h0)]))),
              (-(~^(&$signed(reg1122))))};
          reg1140 <= {reg1129[(4'hb):(2'h2)],
              $unsigned($signed((wire871[(4'hf):(4'hd)] * (~&(8'h9c)))))};
        end
      for (forvar1141 = (1'h0); (forvar1141 < (2'h3)); forvar1141 = (forvar1141 + (1'h1)))
        begin
          for (forvar1142 = (1'h0); (forvar1142 < (1'h0)); forvar1142 = (forvar1142 + (1'h1)))
            begin
              reg1143 <= $unsigned((reg1114 == reg987));
            end
          reg1144 <= (8'h9c);
          reg1145 = (~(8'ha2));
          for (forvar1146 = (1'h0); (forvar1146 < (2'h2)); forvar1146 = (forvar1146 + (1'h1)))
            begin
              reg1147 <= {((~&(!(wire984 ?
                      reg1119 : wire869))) != $unsigned($unsigned((reg879 + reg1129)))),
                  reg1143[(4'ha):(3'h5)]};
              reg1148 <= $signed(((&(((8'hb6) ? wire985 : reg1114) ?
                      (wire1132 ? wire869 : reg1065) : (~(8'h9d)))) ?
                  (-$signed($signed(reg1129))) : ($signed(wire869[(5'h10):(2'h2)]) - forvar1146)));
              reg1149 = reg990[(3'h4):(2'h3)];
              reg1150 <= (8'hba);
            end
        end
      reg1151 = $unsigned(reg1147[(4'hd):(4'hb)]);
      reg1152 = $signed((~|(^$signed((~&(8'h9d))))));
    end
  always
    @(posedge clk) begin
      reg1153 <= forvar874;
      reg1154 = ($signed({wire1108[(4'h9):(4'h9)]}) + $signed(({(forvar991 == reg1069),
              (wire935 ? reg1126 : reg1111)} ?
          {reg1130} : (!$unsigned(wire1062)))));
      reg1155 = $signed($signed(({(8'ha4),
          $signed((8'ha5))} || $unsigned($signed(reg993)))));
      reg1156 <= (reg1124 ? reg1068[(4'hd):(1'h0)] : $unsigned(reg992));
      for (forvar1157 = (1'h0); (forvar1157 < (2'h2)); forvar1157 = (forvar1157 + (1'h1)))
        begin
          reg1158 <= {$signed(reg1069[(3'h7):(1'h0)]),
              ((8'ha4) ?
                  ((~&reg1120[(4'h8):(3'h5)]) ?
                      reg1124 : ($signed(wire1127) ?
                          reg880[(3'h6):(2'h2)] : $unsigned(forvar1157))) : reg1071)};
          reg1159 <= reg1154[(2'h2):(1'h0)];
          reg1160 <= ((wire1073 * {(^~$unsigned(reg1144))}) ?
              forvar1112 : {$unsigned(((~^wire1127) ?
                      $signed(reg1124) : (forvar1157 >> reg1130))),
                  $signed({(reg1148 ? wire1073 : reg1144),
                      $unsigned(wire1132)})});
          reg1161 = $unsigned($signed(reg987[(1'h1):(1'h1)]));
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1074
#( parameter param1106 = {{((~&((8'hba) ? (8'hbe) : (8'ha5))) ? {((8'ha4) ? (8'hae) : (8'ha2)), ((8'hb0) ? (8'h9c) : (8'hb1))} : (((8'ha8) ? (8'h9e) : (8'ha6)) ? {(8'ha8)} : (-(8'ha4))))}, ((((!(8'ha4)) ? {(8'hb9)} : {(8'hb5), (8'hac)}) ? (((8'ha2) ^ (8'ha4)) != (^(7'h42))) : ((~|(8'hac)) > {(8'hae), (8'ha8)})) >> (|((!(7'h44)) + (-(8'ha7)))))}
, parameter param1107 = param1106 )
(y, clk, wire1078, wire1077, wire1076, wire1075);
  output wire [(32'h14e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire1078;
  input wire signed [(2'h2):(1'h0)] wire1077;
  input wire signed [(2'h3):(1'h0)] wire1076;
  input wire [(4'hb):(1'h0)] wire1075;
  wire signed [(5'h10):(1'h0)] wire1105;
  wire signed [(3'h6):(1'h0)] wire1104;
  reg signed [(3'h4):(1'h0)] reg1103 = (1'h0);
  reg [(5'h11):(1'h0)] reg1102 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1101 = (1'h0);
  reg [(4'he):(1'h0)] reg1100 = (1'h0);
  reg [(5'h14):(1'h0)] reg1099 = (1'h0);
  reg [(5'h12):(1'h0)] reg1098 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar1095 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1097 = (1'h0);
  reg [(5'h14):(1'h0)] reg1096 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1095 = (1'h0);
  reg [(5'h15):(1'h0)] reg1094 = (1'h0);
  reg [(2'h3):(1'h0)] reg1093 = (1'h0);
  reg [(3'h7):(1'h0)] reg1092 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1091 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1090 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1089 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1088 = (1'h0);
  reg [(4'hd):(1'h0)] reg1087 = (1'h0);
  reg [(4'hf):(1'h0)] reg1086 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1085 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1084 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1083 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1082 = (1'h0);
  reg [(2'h2):(1'h0)] reg1081 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1080 = (1'h0);
  reg [(2'h2):(1'h0)] reg1079 = (1'h0);
  assign y = {wire1105,
                 wire1104,
                 reg1103,
                 reg1102,
                 forvar1101,
                 reg1100,
                 reg1099,
                 reg1098,
                 forvar1095,
                 reg1097,
                 reg1096,
                 reg1095,
                 reg1094,
                 reg1093,
                 reg1092,
                 reg1091,
                 reg1090,
                 forvar1089,
                 reg1088,
                 reg1087,
                 reg1086,
                 reg1085,
                 forvar1084,
                 reg1083,
                 reg1082,
                 reg1081,
                 forvar1080,
                 reg1079,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1079 = (^wire1075);
      for (forvar1080 = (1'h0); (forvar1080 < (2'h3)); forvar1080 = (forvar1080 + (1'h1)))
        begin
          reg1081 <= wire1076;
          reg1082 <= forvar1080;
        end
      reg1083 <= (({wire1075[(1'h0):(1'h0)]} ?
              ((7'h40) >> ($signed(wire1077) ^~ reg1081)) : (wire1075[(3'h7):(3'h5)] ?
                  wire1077 : wire1077)) ?
          $signed((((~^wire1078) ?
              $unsigned(reg1079) : $unsigned(reg1082)) >>> wire1078)) : ($unsigned($signed(wire1077[(2'h2):(1'h1)])) ?
              reg1079 : {(forvar1080 & $unsigned(wire1078)),
                  $unsigned((wire1077 - forvar1080))}));
    end
  always
    @(posedge clk) begin
      for (forvar1084 = (1'h0); (forvar1084 < (1'h1)); forvar1084 = (forvar1084 + (1'h1)))
        begin
          reg1085 <= $unsigned(((((forvar1080 && (8'ha3)) ?
              $unsigned((8'h9f)) : (reg1081 * forvar1084)) <<< ((~(7'h40)) + reg1081)) * (8'hb5)));
          reg1086 <= (((|(wire1075 ?
              $signed(wire1077) : (&(8'hb0)))) >>> ($signed(((8'ha7) << (8'ha7))) ?
              ($signed(reg1079) < reg1081) : (+(reg1081 ?
                  reg1085 : (8'hab))))) >> wire1077[(1'h1):(1'h0)]);
          reg1087 <= reg1083[(1'h0):(1'h0)];
          reg1088 = (~&{$unsigned(forvar1084)});
          for (forvar1089 = (1'h0); (forvar1089 < (3'h4)); forvar1089 = (forvar1089 + (1'h1)))
            begin
              reg1090 <= ((forvar1089 ?
                  $signed(reg1082[(5'h11):(4'h9)]) : wire1075) >>> ((~|{(reg1088 & forvar1080),
                  (~(8'hb5))}) < reg1085));
              reg1091 = reg1083[(1'h0):(1'h0)];
              reg1092 <= (reg1081 ?
                  (reg1085[(2'h3):(1'h1)] ?
                      ($signed($signed(forvar1080)) ^~ $signed((reg1083 > reg1086))) : $unsigned(reg1086[(4'hb):(3'h4)])) : (($signed({reg1085}) + reg1086[(4'hd):(3'h5)]) ?
                      ((+(forvar1089 | wire1078)) ?
                          $unsigned(reg1087) : reg1082[(3'h5):(3'h5)]) : ((reg1079[(2'h2):(1'h1)] ?
                              $unsigned((8'hb4)) : (~&reg1085)) ?
                          wire1076 : (~reg1081[(2'h2):(1'h0)]))));
            end
        end
      reg1093 <= {$signed(forvar1080),
          (-($signed((reg1081 - (8'h9e))) ?
              ($signed(wire1076) > ((8'hbd) != reg1082)) : reg1092[(3'h5):(2'h3)]))};
      reg1094 <= $signed({(~{(reg1090 && reg1087)})});
      if (($unsigned((($unsigned(reg1086) ?
          reg1086[(4'ha):(3'h6)] : reg1090[(4'ha):(4'h8)]) >>> $signed(reg1081))) ^ (reg1088[(1'h0):(1'h0)] || $unsigned($unsigned((+wire1077))))))
        begin
          reg1095 <= $signed(({(~|(~^wire1077)),
              $signed((reg1086 < (8'hb2)))} != $unsigned($signed($unsigned(reg1091)))));
          reg1096 <= (-({reg1086, reg1083} ?
              $unsigned(((-reg1093) ?
                  (reg1082 < reg1088) : reg1081)) : forvar1084[(2'h3):(1'h1)]));
          reg1097 = $signed(forvar1080[(3'h5):(3'h5)]);
        end
      else
        begin
          for (forvar1095 = (1'h0); (forvar1095 < (1'h0)); forvar1095 = (forvar1095 + (1'h1)))
            begin
              reg1096 <= (8'hba);
              reg1097 <= $unsigned(($signed(reg1079[(1'h1):(1'h0)]) ?
                  $unsigned($signed(reg1085)) : reg1085[(3'h5):(1'h1)]));
              reg1098 <= $signed($unsigned($unsigned((^~reg1086[(3'h7):(1'h1)]))));
              reg1099 <= {(((reg1098 ?
                          ((8'h9f) ?
                              wire1078 : reg1086) : (7'h44)) > (~(reg1093 << reg1083))) ?
                      $signed(($signed(forvar1084) ?
                          reg1087[(2'h2):(2'h2)] : reg1082[(4'hc):(2'h2)])) : (^~reg1082[(4'he):(3'h5)]))};
            end
          reg1100 <= $unsigned((8'ha8));
          for (forvar1101 = (1'h0); (forvar1101 < (2'h2)); forvar1101 = (forvar1101 + (1'h1)))
            begin
              reg1102 <= reg1096[(4'ha):(3'h7)];
            end
        end
      reg1103 <= (reg1093 ?
          reg1090[(4'he):(3'h6)] : $signed($signed($signed(reg1082[(5'h12):(4'h9)]))));
    end
  assign wire1104 = (($unsigned(((reg1092 && reg1094) <= (reg1086 <= reg1099))) && ((~&reg1081[(1'h1):(1'h0)]) ?
                            ($signed(wire1078) ?
                                (-wire1077) : (wire1077 != forvar1084)) : {{reg1090,
                                    reg1083},
                                $unsigned(reg1088)})) ?
                        reg1083 : (|({$unsigned(wire1078),
                            (forvar1089 + wire1075)} && reg1092)));
  assign wire1105 = {$signed(wire1077)};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module994  (y, clk, wire999, wire998, wire997, wire996, wire995);
  output wire [(32'h2d3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h7):(1'h0)] wire999;
  input wire [(3'h7):(1'h0)] wire998;
  input wire signed [(3'h6):(1'h0)] wire997;
  input wire signed [(4'hf):(1'h0)] wire996;
  input wire signed [(5'h12):(1'h0)] wire995;
  reg [(3'h7):(1'h0)] reg1061 = (1'h0);
  reg [(4'hc):(1'h0)] reg1060 = (1'h0);
  reg [(4'ha):(1'h0)] reg1059 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1058 = (1'h0);
  wire [(4'hb):(1'h0)] wire1057;
  reg [(3'h7):(1'h0)] reg1056 = (1'h0);
  reg [(3'h6):(1'h0)] reg1055 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1054 = (1'h0);
  reg [(5'h10):(1'h0)] reg1053 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1052 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1050 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1051 = (1'h0);
  reg [(4'hb):(1'h0)] reg1050 = (1'h0);
  reg [(4'hf):(1'h0)] reg1049 = (1'h0);
  reg [(3'h5):(1'h0)] reg1048 = (1'h0);
  reg [(5'h10):(1'h0)] reg1047 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1046 = (1'h0);
  reg [(2'h3):(1'h0)] reg1045 = (1'h0);
  reg [(4'he):(1'h0)] forvar1044 = (1'h0);
  reg [(4'he):(1'h0)] reg1043 = (1'h0);
  reg [(5'h14):(1'h0)] reg1042 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1041 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1040 = (1'h0);
  reg [(3'h5):(1'h0)] reg1039 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1038 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1037 = (1'h0);
  reg [(3'h4):(1'h0)] reg1036 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1035 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire1034;
  reg [(2'h3):(1'h0)] reg1033 = (1'h0);
  reg [(4'hd):(1'h0)] reg1032 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1031 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1030 = (1'h0);
  reg [(4'ha):(1'h0)] reg1029 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1028 = (1'h0);
  reg [(3'h4):(1'h0)] reg1027 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire1026;
  reg [(3'h7):(1'h0)] reg1025 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1024 = (1'h0);
  wire [(5'h10):(1'h0)] wire1023;
  wire [(2'h2):(1'h0)] wire1022;
  reg signed [(4'hb):(1'h0)] reg1021 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1020 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1019 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire1018;
  reg [(5'h11):(1'h0)] reg1017 = (1'h0);
  reg [(2'h2):(1'h0)] reg1016 = (1'h0);
  reg [(5'h12):(1'h0)] reg1015 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire1014;
  wire signed [(3'h6):(1'h0)] wire1013;
  reg signed [(5'h12):(1'h0)] reg1012 = (1'h0);
  reg [(4'h8):(1'h0)] reg1011 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire1010;
  reg [(5'h11):(1'h0)] reg1009 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1003 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1002 = (1'h0);
  reg [(5'h10):(1'h0)] reg1008 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1007 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1006 = (1'h0);
  reg [(4'hd):(1'h0)] reg1005 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1004 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1003 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1002 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1001 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1000 = (1'h0);
  assign y = {reg1061,
                 reg1060,
                 reg1059,
                 reg1058,
                 wire1057,
                 reg1056,
                 reg1055,
                 reg1054,
                 reg1053,
                 reg1052,
                 forvar1050,
                 reg1051,
                 reg1050,
                 reg1049,
                 reg1048,
                 reg1047,
                 reg1046,
                 reg1045,
                 forvar1044,
                 reg1043,
                 reg1042,
                 reg1041,
                 reg1040,
                 reg1039,
                 reg1038,
                 forvar1037,
                 reg1036,
                 forvar1035,
                 wire1034,
                 reg1033,
                 reg1032,
                 reg1031,
                 reg1030,
                 reg1029,
                 forvar1028,
                 reg1027,
                 wire1026,
                 reg1025,
                 reg1024,
                 wire1023,
                 wire1022,
                 reg1021,
                 reg1020,
                 reg1019,
                 wire1018,
                 reg1017,
                 reg1016,
                 reg1015,
                 wire1014,
                 wire1013,
                 reg1012,
                 reg1011,
                 wire1010,
                 reg1009,
                 reg1003,
                 forvar1002,
                 reg1008,
                 reg1007,
                 reg1006,
                 reg1005,
                 reg1004,
                 forvar1003,
                 reg1002,
                 reg1001,
                 reg1000,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ((-($unsigned((^~wire996)) ?
          (wire999[(1'h0):(1'h0)] ?
              ((wire996 | wire998) ?
                  {wire995} : (wire997 == wire995)) : $unsigned((wire995 ?
                  (8'haf) : wire998))) : wire999[(1'h0):(1'h0)])))
        begin
          reg1000 <= wire998[(1'h1):(1'h1)];
          reg1001 <= $unsigned((+wire995));
          reg1002 <= reg1001[(4'hb):(1'h0)];
          for (forvar1003 = (1'h0); (forvar1003 < (1'h1)); forvar1003 = (forvar1003 + (1'h1)))
            begin
              reg1004 <= (7'h41);
              reg1005 <= wire998[(1'h1):(1'h1)];
              reg1006 = ((wire997[(3'h5):(1'h0)] ?
                  $unsigned($unsigned(((8'ha5) == wire995))) : (^((|wire997) >>> wire999))) >> (forvar1003 ?
                  reg1002[(3'h6):(2'h2)] : {(|$signed(reg1004)),
                      $unsigned(((8'hbb) ^~ reg1000))}));
              reg1007 = $unsigned(((~&($signed((8'hb2)) ?
                  reg1000 : $unsigned((8'hb1)))) > $signed($signed((8'hba)))));
            end
          reg1008 = ($unsigned(wire999) ? wire995 : reg1001[(4'h9):(2'h3)]);
        end
      else
        begin
          reg1000 <= $unsigned($unsigned($signed(wire997)));
          reg1001 <= (~|$signed((reg1002[(1'h1):(1'h0)] > ((reg1004 ?
              reg1007 : reg1006) | reg1001[(3'h5):(3'h4)]))));
          for (forvar1002 = (1'h0); (forvar1002 < (2'h2)); forvar1002 = (forvar1002 + (1'h1)))
            begin
              reg1003 <= wire996;
              reg1004 <= (~|($unsigned($unsigned((^reg1006))) > $signed(forvar1002[(3'h4):(3'h4)])));
              reg1005 <= reg1007[(4'h9):(4'h9)];
            end
          reg1006 <= (8'ha7);
        end
    end
  always
    @(posedge clk) begin
      reg1009 <= (&((!((|reg1002) == (!reg1000))) != $signed($unsigned((+forvar1002)))));
    end
  assign wire1010 = ((wire998 <= reg1007[(3'h5):(1'h1)]) > ($signed(reg1007[(3'h4):(3'h4)]) ?
                        $unsigned({(^reg1006)}) : (($signed((8'hbe)) <<< (&reg1007)) ?
                            forvar1003 : wire998)));
  always
    @(posedge clk) begin
      reg1011 <= $signed(wire1010[(2'h3):(2'h3)]);
      reg1012 <= {(reg1007[(5'h13):(4'hb)] ?
              forvar1003[(2'h3):(2'h2)] : reg1005),
          $unsigned(wire998)};
    end
  assign wire1013 = (reg1012 ?
                        reg1004[(2'h3):(1'h1)] : ($unsigned($signed($unsigned(wire997))) ?
                            (!wire999) : ($signed({(7'h42)}) != reg1012[(4'h9):(2'h3)])));
  assign wire1014 = $signed((reg1000 >>> forvar1002[(2'h3):(1'h0)]));
  always
    @(posedge clk) begin
      reg1015 = $unsigned({(wire997 ? wire998 : reg1004),
          ($unsigned(wire1013[(3'h6):(2'h2)]) <<< $unsigned((wire996 | wire997)))});
    end
  always
    @(posedge clk) begin
      reg1016 <= reg1000;
      reg1017 = $unsigned($unsigned(reg1006[(1'h1):(1'h1)]));
    end
  assign wire1018 = $signed((8'hb2));
  always
    @(posedge clk) begin
      reg1019 = ((~&({(reg1002 ?
              (8'hb6) : reg1002)} ^~ {$unsigned(forvar1003)})) >>> forvar1002);
      reg1020 = $signed(reg1002);
      reg1021 = wire997;
    end
  assign wire1022 = wire995;
  assign wire1023 = {{reg1019},
                        $signed($unsigned($unsigned($unsigned((8'hb2)))))};
  always
    @(posedge clk) begin
      reg1024 = (wire1023 ?
          (^reg1016) : $unsigned((wire997[(3'h6):(2'h2)] <<< (wire995[(3'h4):(2'h3)] ?
              (reg1003 & reg1005) : $unsigned(reg1008)))));
      reg1025 = (($signed((8'hbc)) >= $signed(({reg1015} || $unsigned((8'h9d))))) ?
          wire1013 : ((((8'hb4) >>> (~^reg1008)) >= (8'ha6)) * $signed({{reg1001,
                  reg1004}})));
    end
  assign wire1026 = reg1009[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      reg1027 <= $unsigned((-reg1017));
      for (forvar1028 = (1'h0); (forvar1028 < (2'h3)); forvar1028 = (forvar1028 + (1'h1)))
        begin
          reg1029 = {wire1018};
          reg1030 = $unsigned(reg1021);
          reg1031 <= forvar1003;
        end
      reg1032 <= reg1030;
      reg1033 <= ($unsigned($signed($unsigned((&(8'ha8))))) | $signed(reg1009));
    end
  assign wire1034 = {$signed($unsigned($unsigned((+(8'hbd))))), wire998};
  always
    @(posedge clk) begin
      for (forvar1035 = (1'h0); (forvar1035 < (1'h1)); forvar1035 = (forvar1035 + (1'h1)))
        begin
          reg1036 <= (reg1021 > (reg1021[(3'h7):(2'h3)] ?
              $unsigned($unsigned((|(8'hbb)))) : (^~(|$signed(reg1005)))));
          for (forvar1037 = (1'h0); (forvar1037 < (3'h4)); forvar1037 = (forvar1037 + (1'h1)))
            begin
              reg1038 <= $signed((8'ha7));
            end
          reg1039 <= {$signed($unsigned($signed($signed(reg1038)))),
              (reg1015 != (^~((!reg1012) >> {forvar1002, reg1032})))};
          reg1040 <= {{{(-reg1002[(4'he):(3'h7)]), (~^((8'hae) > reg1029))}}};
          reg1041 <= $unsigned(reg1029);
        end
      reg1042 <= reg1024[(4'h8):(1'h0)];
      if (forvar1002)
        begin
          reg1043 <= ((wire998[(2'h3):(2'h3)] ?
              wire997[(2'h3):(1'h1)] : $unsigned(wire1026)) * reg1024);
          for (forvar1044 = (1'h0); (forvar1044 < (2'h2)); forvar1044 = (forvar1044 + (1'h1)))
            begin
              reg1045 <= forvar1003;
              reg1046 <= ({$unsigned((8'h9d))} ?
                  ($signed(((forvar1002 ? (8'ha1) : wire1026) ?
                      $unsigned(reg1011) : reg1040)) | (forvar1002 ?
                      ($unsigned(wire1010) > (~&reg1019)) : $unsigned({forvar1037}))) : reg1027);
              reg1047 = ((+((~&(8'hba)) ?
                  ($unsigned(wire997) - wire1010[(3'h4):(1'h0)]) : ($signed(reg1032) ?
                      reg1032 : $signed((8'ha7))))) & (({$signed(reg1046)} < reg1009) < $unsigned(reg1001)));
              reg1048 <= reg1024;
              reg1049 <= $unsigned((~^(~^{reg1031[(4'hc):(4'h8)]})));
            end
          reg1050 <= (|{wire997, $unsigned($unsigned($unsigned(reg1006)))});
          reg1051 <= {((~^((~|wire996) ?
                  (reg1020 ?
                      reg1002 : reg1001) : (^~forvar1003))) ^~ $signed(((reg1020 >>> wire1023) ?
                  reg1016[(1'h1):(1'h1)] : {reg1029})))};
        end
      else
        begin
          reg1043 = $signed((&((reg1045[(2'h2):(1'h0)] << $unsigned(reg1009)) ?
              reg1021 : ($unsigned((8'hbd)) ?
                  wire995[(4'h9):(2'h2)] : {(8'h9c)}))));
          for (forvar1044 = (1'h0); (forvar1044 < (2'h2)); forvar1044 = (forvar1044 + (1'h1)))
            begin
              reg1045 = (7'h43);
              reg1046 = $unsigned(forvar1037[(2'h2):(1'h0)]);
              reg1047 = (~&forvar1003);
              reg1048 <= (~^reg1045[(2'h2):(2'h2)]);
            end
          reg1049 <= (({$unsigned($unsigned(reg1005))} ?
              {reg1007[(5'h11):(1'h1)]} : reg1024) > ((reg1027[(2'h2):(2'h2)] >= reg1041[(1'h1):(1'h1)]) ?
              (7'h40) : reg1031[(3'h7):(3'h5)]));
          for (forvar1050 = (1'h0); (forvar1050 < (2'h3)); forvar1050 = (forvar1050 + (1'h1)))
            begin
              reg1051 <= (8'hb2);
              reg1052 = {(8'ha5)};
              reg1053 = (&$signed((($signed(reg1024) || forvar1003[(3'h4):(3'h4)]) ?
                  $unsigned((~(8'ha9))) : reg1040[(1'h0):(1'h0)])));
              reg1054 <= ((($signed((reg1016 <= reg1012)) + (reg1047 ^ $unsigned(forvar1028))) ~^ $unsigned((8'hb5))) ?
                  {forvar1002[(4'h9):(3'h6)],
                      $signed({(wire1018 + (7'h40))})} : (8'hb8));
            end
          reg1055 <= {{$signed(((reg1019 != forvar1035) ^~ ((7'h40) >= reg1020))),
                  forvar1003[(2'h2):(2'h2)]}};
        end
      reg1056 <= ({reg1033, (~|$unsigned(reg1003))} ?
          $unsigned((~wire1022)) : reg1050);
    end
  assign wire1057 = (8'hb8);
  always
    @(posedge clk) begin
      reg1058 <= (!(~&$signed(((~^reg1008) > $unsigned((8'hb3))))));
      reg1059 <= (^~((^((reg1009 != reg1051) >= $signed((7'h43)))) ?
          reg1036[(2'h2):(2'h2)] : ((^((8'ha9) <= wire1026)) | (~|{(8'ha4),
              reg1041}))));
      reg1060 <= ((((!(reg1032 <<< reg1031)) >= reg1003) | reg1004) ?
          $signed($unsigned(($signed(forvar1028) + (~|reg1002)))) : reg1011[(1'h1):(1'h0)]);
      reg1061 = $unsigned($signed(({$unsigned(forvar1035)} ?
          $signed(((8'hb0) + reg1049)) : ($signed(wire995) ^ (reg1036 + reg1038)))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module937
#( parameter param980 = ((&(8'had)) < (((~&(~^(8'hb4))) ? (^~(~|(8'hb4))) : (((8'hbf) ? (8'hbb) : (8'ha0)) ^~ ((8'hae) != (8'hae)))) ? (((~^(8'hb8)) ? ((7'h44) != (8'hb6)) : (8'hbc)) ? (!{(8'haa), (8'hb3)}) : (-((8'ha7) ^ (8'ha1)))) : ({((8'haf) ~^ (8'hac)), ((8'hb5) ? (8'hb5) : (8'hb8))} ? (-{(8'hb3)}) : (&(+(8'h9c))))))
, parameter param981 = param980 )
(y, clk, wire941, wire940, wire939, wire938);
  output wire [(32'h1aa):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire941;
  input wire [(4'hf):(1'h0)] wire940;
  input wire [(5'h13):(1'h0)] wire939;
  input wire [(5'h12):(1'h0)] wire938;
  wire signed [(4'h8):(1'h0)] wire979;
  wire signed [(4'h8):(1'h0)] wire978;
  reg signed [(4'h9):(1'h0)] reg977 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg976 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg975 = (1'h0);
  reg signed [(4'he):(1'h0)] reg972 = (1'h0);
  reg [(5'h11):(1'h0)] reg974 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg973 = (1'h0);
  reg [(4'hf):(1'h0)] forvar972 = (1'h0);
  reg [(4'h9):(1'h0)] reg971 = (1'h0);
  reg [(4'hd):(1'h0)] reg970 = (1'h0);
  reg [(3'h7):(1'h0)] reg969 = (1'h0);
  reg [(4'h9):(1'h0)] reg968 = (1'h0);
  wire [(3'h4):(1'h0)] wire967;
  wire [(3'h7):(1'h0)] wire966;
  wire signed [(3'h4):(1'h0)] wire965;
  reg signed [(4'hc):(1'h0)] reg964 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg963 = (1'h0);
  reg [(3'h6):(1'h0)] reg962 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg961 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg960 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar959 = (1'h0);
  reg [(3'h4):(1'h0)] reg958 = (1'h0);
  reg [(4'h8):(1'h0)] reg957 = (1'h0);
  wire [(3'h4):(1'h0)] wire956;
  wire signed [(2'h2):(1'h0)] wire955;
  wire [(3'h5):(1'h0)] wire954;
  reg signed [(5'h12):(1'h0)] reg953 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg952 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg951 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg950 = (1'h0);
  reg [(5'h14):(1'h0)] forvar949 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg948 = (1'h0);
  wire [(5'h15):(1'h0)] wire947;
  reg [(4'hd):(1'h0)] reg946 = (1'h0);
  reg [(4'h8):(1'h0)] reg945 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg944 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar943 = (1'h0);
  reg [(4'hf):(1'h0)] reg942 = (1'h0);
  assign y = {wire979,
                 wire978,
                 reg977,
                 reg976,
                 reg975,
                 reg972,
                 reg974,
                 reg973,
                 forvar972,
                 reg971,
                 reg970,
                 reg969,
                 reg968,
                 wire967,
                 wire966,
                 wire965,
                 reg964,
                 reg963,
                 reg962,
                 reg961,
                 reg960,
                 forvar959,
                 reg958,
                 reg957,
                 wire956,
                 wire955,
                 wire954,
                 reg953,
                 reg952,
                 reg951,
                 reg950,
                 forvar949,
                 reg948,
                 wire947,
                 reg946,
                 reg945,
                 reg944,
                 forvar943,
                 reg942,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg942 <= wire941;
      for (forvar943 = (1'h0); (forvar943 < (2'h3)); forvar943 = (forvar943 + (1'h1)))
        begin
          reg944 <= $unsigned($unsigned((+((forvar943 < wire940) ~^ (!wire938)))));
        end
      reg945 <= wire938[(5'h10):(4'hb)];
      reg946 = reg944[(3'h5):(2'h3)];
    end
  assign wire947 = wire940[(4'h9):(1'h0)];
  always
    @(posedge clk) begin
      reg948 <= ({(-wire947[(3'h5):(2'h3)])} ~^ ($unsigned((reg944[(3'h7):(1'h0)] ?
          wire947[(3'h4):(3'h4)] : $signed(wire947))) != (~^((forvar943 != wire947) <<< wire939))));
      for (forvar949 = (1'h0); (forvar949 < (1'h1)); forvar949 = (forvar949 + (1'h1)))
        begin
          reg950 <= ($signed(($signed((reg944 ? forvar943 : wire939)) ?
              ({forvar949, (8'hab)} + reg942) : wire938)) >>> reg944);
          reg951 = ($unsigned(wire941) ?
              (~&{(8'ha0)}) : (reg948[(1'h1):(1'h1)] ?
                  ({(wire941 - reg948)} ^ reg946) : wire947));
        end
      reg952 <= (~&(forvar943[(5'h11):(4'h8)] ~^ {($signed(reg942) > $unsigned(forvar949))}));
      reg953 <= (((reg944[(3'h4):(1'h0)] ~^ $signed(reg942)) ?
          (reg952 ?
              (reg951 >>> wire939) : ($signed((8'haa)) ~^ (^~reg946))) : reg942[(3'h6):(1'h0)]) != $signed(((8'hbb) ?
          (^~reg952[(4'h9):(1'h0)]) : {$signed(reg948)})));
    end
  assign wire954 = $signed({(^(~^(&reg948))), (reg952 >> forvar943)});
  assign wire955 = reg944[(1'h0):(1'h0)];
  assign wire956 = $unsigned(wire954[(1'h1):(1'h0)]);
  always
    @(posedge clk) begin
      reg957 <= wire941;
      reg958 <= (wire956 & ((^~$unsigned((+reg948))) ?
          ({{wire938, reg957}} ?
              $signed(reg952[(2'h3):(2'h2)]) : (8'hb9)) : wire938[(1'h1):(1'h0)]));
      for (forvar959 = (1'h0); (forvar959 < (3'h4)); forvar959 = (forvar959 + (1'h1)))
        begin
          reg960 = (reg948[(3'h4):(1'h1)] ?
              {(($unsigned(reg948) == reg957) ?
                      $unsigned(wire940) : (!forvar949)),
                  ((7'h44) + wire938[(1'h1):(1'h1)])} : (|reg944[(1'h0):(1'h0)]));
          reg961 <= wire939;
          reg962 <= $signed($signed((forvar949[(4'h8):(3'h7)] < {$unsigned((8'hb9))})));
        end
      reg963 = forvar943[(4'h8):(1'h1)];
      reg964 = ((+reg957) ?
          $unsigned($signed((|(~reg953)))) : $signed((~^(~^reg960))));
    end
  assign wire965 = wire938[(5'h10):(3'h6)];
  assign wire966 = reg964;
  assign wire967 = reg952[(3'h6):(3'h6)];
  always
    @(posedge clk) begin
      reg968 = $signed(reg957[(2'h3):(2'h2)]);
      reg969 <= ((($unsigned((8'hb9)) >>> (((8'hbd) ? wire938 : reg963) ?
              {reg948, wire941} : reg952)) ?
          (~reg961[(4'hd):(4'h9)]) : (wire954[(1'h0):(1'h0)] ?
              wire941[(4'hc):(2'h3)] : $signed($signed(wire954)))) | (|wire941));
      reg970 <= ($unsigned(($unsigned((forvar949 >> reg946)) >> (~|$signed(wire947)))) ?
          {(8'ha9),
              $signed(reg961)} : $signed($signed($unsigned((reg951 != (8'h9e))))));
      reg971 <= $signed(reg952[(5'h14):(4'h9)]);
    end
  always
    @(posedge clk) begin
      if ($unsigned((+($unsigned($unsigned(wire947)) ?
          ($unsigned(reg968) ?
              (reg951 | wire955) : $unsigned(reg960)) : (^$unsigned(wire954))))))
        begin
          for (forvar972 = (1'h0); (forvar972 < (2'h2)); forvar972 = (forvar972 + (1'h1)))
            begin
              reg973 <= reg952[(4'hd):(4'h8)];
            end
          reg974 <= (wire955[(2'h2):(1'h0)] ?
              $signed(wire939) : $unsigned(($unsigned((!reg970)) ?
                  ((~(7'h44)) ?
                      reg951[(2'h2):(2'h2)] : wire954) : {$unsigned(forvar959)})));
        end
      else
        begin
          reg972 <= (forvar943 ?
              $unsigned({(reg964 << (reg944 ?
                      wire941 : (8'hb1)))}) : wire938[(4'h9):(3'h6)]);
          reg973 <= (^reg946);
        end
      reg975 = ((reg968 ? reg952 : forvar949) ?
          (~&reg973[(3'h7):(1'h0)]) : ((((reg968 ?
                  wire965 : wire938) - $signed((8'hb6))) ?
              $signed($unsigned((8'hbd))) : (^{(7'h42), reg962})) << ((8'hbf) ?
              ((8'h9e) ?
                  (reg953 ?
                      reg972 : reg969) : (~|reg962)) : $signed($unsigned(reg970)))));
      reg976 = wire941[(4'h8):(3'h5)];
      reg977 <= (($signed((wire940[(3'h6):(3'h6)] ?
              reg961[(5'h11):(4'ha)] : (|reg975))) ?
          reg945 : $unsigned((~|reg948))) <<< reg972);
    end
  assign wire978 = (wire967 ?
                       reg974[(5'h10):(5'h10)] : ((8'h9c) ?
                           ((!wire940) ?
                               ((~&wire941) ?
                                   $unsigned(forvar959) : (+wire966)) : $signed($signed(reg963))) : $unsigned(wire967)));
  assign wire979 = ({(($unsigned(reg960) ?
                                   reg975[(1'h1):(1'h1)] : $signed(reg964)) ?
                               forvar972 : {forvar959, reg976[(2'h3):(2'h2)]}),
                           $signed((((8'haa) ? reg963 : reg957) ?
                               (8'ha7) : (reg948 || reg950)))} ?
                       $signed(reg950[(3'h6):(3'h6)]) : reg969);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module881
#(parameter param934 = (~(8'hbb)))
(y, clk, wire886, wire885, wire884, wire883, wire882);
  output wire [(32'h256):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h7):(1'h0)] wire886;
  input wire [(2'h3):(1'h0)] wire885;
  input wire signed [(4'hc):(1'h0)] wire884;
  input wire signed [(5'h12):(1'h0)] wire883;
  input wire [(4'h8):(1'h0)] wire882;
  wire [(5'h15):(1'h0)] wire933;
  reg [(5'h14):(1'h0)] reg932 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg931 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg930 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg929 = (1'h0);
  reg [(3'h7):(1'h0)] reg928 = (1'h0);
  reg [(4'ha):(1'h0)] reg927 = (1'h0);
  reg signed [(4'he):(1'h0)] reg926 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg925 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg924 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg923 = (1'h0);
  reg [(4'h8):(1'h0)] reg922 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg921 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire920;
  reg [(5'h10):(1'h0)] reg919 = (1'h0);
  reg [(4'h8):(1'h0)] reg918 = (1'h0);
  reg [(5'h13):(1'h0)] reg917 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg916 = (1'h0);
  reg [(3'h6):(1'h0)] forvar915 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg914 = (1'h0);
  reg [(4'h9):(1'h0)] reg913 = (1'h0);
  reg [(2'h3):(1'h0)] reg912 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg911 = (1'h0);
  reg [(3'h4):(1'h0)] reg910 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg909 = (1'h0);
  reg [(5'h10):(1'h0)] forvar908 = (1'h0);
  wire [(3'h6):(1'h0)] wire907;
  wire [(4'hb):(1'h0)] wire906;
  wire signed [(4'hb):(1'h0)] wire905;
  reg signed [(4'hd):(1'h0)] reg904 = (1'h0);
  reg [(4'h8):(1'h0)] reg903 = (1'h0);
  reg [(4'hd):(1'h0)] reg902 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg901 = (1'h0);
  reg signed [(4'he):(1'h0)] reg900 = (1'h0);
  reg [(5'h11):(1'h0)] reg899 = (1'h0);
  reg [(4'he):(1'h0)] reg898 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg897 = (1'h0);
  reg [(2'h3):(1'h0)] reg896 = (1'h0);
  reg [(4'ha):(1'h0)] reg895 = (1'h0);
  reg [(4'h9):(1'h0)] reg894 = (1'h0);
  reg [(4'hd):(1'h0)] forvar893 = (1'h0);
  reg [(4'h9):(1'h0)] forvar892 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg891 = (1'h0);
  reg [(3'h5):(1'h0)] reg890 = (1'h0);
  reg [(4'hf):(1'h0)] reg889 = (1'h0);
  reg [(4'hb):(1'h0)] reg888 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar887 = (1'h0);
  assign y = {wire933,
                 reg932,
                 reg931,
                 reg930,
                 reg929,
                 reg928,
                 reg927,
                 reg926,
                 reg925,
                 reg924,
                 reg923,
                 reg922,
                 reg921,
                 wire920,
                 reg919,
                 reg918,
                 reg917,
                 reg916,
                 forvar915,
                 reg914,
                 reg913,
                 reg912,
                 reg911,
                 reg910,
                 reg909,
                 forvar908,
                 wire907,
                 wire906,
                 wire905,
                 reg904,
                 reg903,
                 reg902,
                 reg901,
                 reg900,
                 reg899,
                 reg898,
                 reg897,
                 reg896,
                 reg895,
                 reg894,
                 forvar893,
                 forvar892,
                 reg891,
                 reg890,
                 reg889,
                 reg888,
                 forvar887,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar887 = (1'h0); (forvar887 < (1'h0)); forvar887 = (forvar887 + (1'h1)))
        begin
          reg888 <= (~&wire885);
          reg889 <= (wire885[(2'h3):(2'h3)] ?
              ((~^(&$unsigned(forvar887))) ?
                  $unsigned(({wire885,
                      wire883} ^ $unsigned(forvar887))) : ($signed(wire882[(3'h6):(3'h5)]) ^~ wire884)) : $signed({{(|wire885),
                      ((8'hb6) ? wire884 : forvar887)}}));
          reg890 <= $signed(wire886[(2'h3):(1'h0)]);
        end
      reg891 = (-{$unsigned(($signed(reg888) && $unsigned((8'ha2)))),
          $unsigned($unsigned({reg888}))});
      for (forvar892 = (1'h0); (forvar892 < (1'h0)); forvar892 = (forvar892 + (1'h1)))
        begin
          for (forvar893 = (1'h0); (forvar893 < (3'h4)); forvar893 = (forvar893 + (1'h1)))
            begin
              reg894 <= (~&(+$signed({{forvar893, (8'hab)}, wire882})));
              reg895 = (+({(~^(reg889 | reg894)),
                  wire886[(3'h5):(2'h3)]} - (forvar892 ^ wire883[(4'he):(3'h4)])));
              reg896 <= {{$signed(((wire885 ?
                          (8'hb4) : forvar893) * wire886[(1'h0):(1'h0)])),
                      (|(8'hbd))},
                  forvar893};
              reg897 <= (((+$unsigned((|forvar893))) >= $unsigned(($signed(reg894) - (-wire882)))) ?
                  wire886 : reg889[(4'ha):(1'h1)]);
              reg898 <= reg894;
            end
          reg899 = (reg897 ~^ $unsigned(wire884));
          reg900 = $signed(wire884[(3'h7):(2'h2)]);
          reg901 <= reg897;
          reg902 <= (~{(+($unsigned(reg898) ?
                  $unsigned(reg891) : forvar887[(5'h15):(1'h0)])),
              forvar892});
        end
      reg903 <= wire885;
      reg904 = {reg901[(5'h12):(4'hf)]};
    end
  assign wire905 = $unsigned($signed({$signed((wire886 ? reg897 : (8'had)))}));
  assign wire906 = ($unsigned((8'h9e)) ?
                       wire886[(1'h1):(1'h1)] : (($unsigned($signed(forvar887)) <= forvar887) << (reg894[(1'h0):(1'h0)] ?
                           $unsigned($signed(reg889)) : forvar892)));
  assign wire907 = reg897;
  always
    @(posedge clk) begin
      for (forvar908 = (1'h0); (forvar908 < (1'h1)); forvar908 = (forvar908 + (1'h1)))
        begin
          reg909 = (wire905[(3'h4):(1'h0)] ?
              (($signed({reg894, reg891}) + (wire883[(4'hd):(2'h3)] ?
                      {wire884} : {reg903})) ?
                  ((reg897[(1'h1):(1'h0)] ?
                      {reg904} : ((7'h41) ?
                          forvar908 : reg891)) & ((~forvar887) - wire907)) : (~&reg888)) : ((~&$signed($unsigned(reg890))) < ((^reg894[(1'h1):(1'h0)]) ^ reg902[(4'hb):(3'h7)])));
        end
      reg910 = ($signed(reg909) <= $unsigned(wire886[(3'h7):(3'h7)]));
      reg911 = (^~forvar908);
      reg912 <= wire883;
      reg913 = $signed((reg896 && $unsigned(wire885[(2'h3):(2'h3)])));
    end
  always
    @(posedge clk) begin
      reg914 = reg895;
      for (forvar915 = (1'h0); (forvar915 < (1'h0)); forvar915 = (forvar915 + (1'h1)))
        begin
          reg916 <= reg911;
        end
      reg917 <= wire907[(3'h4):(1'h0)];
      reg918 <= (reg912 ?
          (8'hba) : ($signed((8'hb8)) <= reg917[(3'h5):(1'h1)]));
      reg919 <= (~&wire886);
    end
  assign wire920 = {reg911, wire883[(2'h2):(1'h1)]};
  always
    @(posedge clk) begin
      reg921 <= reg916;
      reg922 = (~reg921[(4'hb):(4'hb)]);
      reg923 <= $signed(reg909[(1'h1):(1'h1)]);
    end
  always
    @(posedge clk) begin
      reg924 <= (reg888[(4'h8):(3'h6)] ?
          $unsigned({reg923,
              forvar893[(3'h7):(3'h4)]}) : (^~reg918[(4'h8):(4'h8)]));
      reg925 <= wire905[(3'h7):(3'h5)];
    end
  always
    @(posedge clk) begin
      if ((+wire885[(1'h0):(1'h0)]))
        begin
          reg926 <= (^~{(~&($signed(reg900) ? $unsigned(reg911) : {wire883}))});
          reg927 = {reg900};
          reg928 = $signed(reg900[(4'h9):(3'h7)]);
        end
      else
        begin
          reg926 = reg921;
        end
      reg929 <= $unsigned(reg898);
      reg930 <= {reg912[(1'h1):(1'h0)], $unsigned(reg903)};
      reg931 <= (~&$unsigned(($signed($unsigned(reg916)) >= ((~(8'hb9)) >>> (~&(8'hbe))))));
      reg932 <= forvar887;
    end
  assign wire933 = $signed(reg900);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1248  (y, clk, wire1252, wire1251, wire1250, wire1249);
  output wire [(32'h1fa):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire1252;
  input wire signed [(4'hc):(1'h0)] wire1251;
  input wire signed [(5'h14):(1'h0)] wire1250;
  input wire signed [(4'he):(1'h0)] wire1249;
  wire signed [(4'hd):(1'h0)] wire1301;
  reg [(4'ha):(1'h0)] reg1300 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1299 = (1'h0);
  wire [(4'h9):(1'h0)] wire1298;
  wire signed [(4'ha):(1'h0)] wire1297;
  reg [(4'ha):(1'h0)] reg1296 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1295 = (1'h0);
  reg [(4'hb):(1'h0)] reg1294 = (1'h0);
  reg [(3'h5):(1'h0)] reg1293 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1292 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire1291;
  reg [(4'hb):(1'h0)] reg1290 = (1'h0);
  reg [(3'h5):(1'h0)] reg1289 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1288 = (1'h0);
  reg [(3'h5):(1'h0)] reg1287 = (1'h0);
  wire [(5'h11):(1'h0)] wire1286;
  reg signed [(3'h6):(1'h0)] reg1285 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1284 = (1'h0);
  reg [(2'h3):(1'h0)] reg1283 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1282 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1281 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1280 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1279 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1278 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1277 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1276 = (1'h0);
  reg [(3'h6):(1'h0)] reg1275 = (1'h0);
  reg [(3'h7):(1'h0)] reg1274 = (1'h0);
  reg [(5'h15):(1'h0)] reg1273 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire1272;
  reg signed [(4'hb):(1'h0)] reg1271 = (1'h0);
  reg [(5'h10):(1'h0)] reg1270 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1269 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1268 = (1'h0);
  reg [(4'h9):(1'h0)] reg1267 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1266 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1265 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire1264;
  wire signed [(5'h11):(1'h0)] wire1263;
  reg signed [(5'h14):(1'h0)] reg1262 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1261 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1260 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1259 = (1'h0);
  reg [(5'h10):(1'h0)] reg1258 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire1257;
  reg [(4'h9):(1'h0)] reg1256 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1255 = (1'h0);
  reg [(4'hb):(1'h0)] reg1254 = (1'h0);
  reg [(2'h3):(1'h0)] reg1253 = (1'h0);
  assign y = {wire1301,
                 reg1300,
                 reg1299,
                 wire1298,
                 wire1297,
                 reg1296,
                 reg1295,
                 reg1294,
                 reg1293,
                 reg1292,
                 wire1291,
                 reg1290,
                 reg1289,
                 forvar1288,
                 reg1287,
                 wire1286,
                 reg1285,
                 reg1284,
                 reg1283,
                 reg1282,
                 reg1281,
                 reg1280,
                 reg1279,
                 reg1278,
                 forvar1277,
                 forvar1276,
                 reg1275,
                 reg1274,
                 reg1273,
                 wire1272,
                 reg1271,
                 reg1270,
                 reg1269,
                 reg1268,
                 reg1267,
                 reg1266,
                 forvar1265,
                 wire1264,
                 wire1263,
                 reg1262,
                 reg1261,
                 reg1260,
                 forvar1259,
                 reg1258,
                 wire1257,
                 reg1256,
                 reg1255,
                 reg1254,
                 reg1253,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1253 <= (+wire1251[(3'h6):(1'h1)]);
      reg1254 <= (~^{$unsigned((wire1251 ?
              (wire1252 | (7'h41)) : $unsigned(wire1249))),
          $unsigned((^(wire1252 ? wire1250 : (7'h43))))});
      reg1255 <= ({wire1249[(2'h3):(2'h3)]} <= reg1253);
      reg1256 <= $signed((wire1250[(1'h0):(1'h0)] ?
          reg1255[(4'hc):(3'h7)] : {wire1249[(3'h4):(2'h2)]}));
    end
  assign wire1257 = (&wire1251);
  always
    @(posedge clk) begin
      reg1258 <= ($unsigned((((wire1249 ? reg1253 : reg1256) ?
              reg1254[(3'h6):(3'h6)] : (reg1253 ?
                  wire1249 : (8'hb8))) == ((wire1250 < (8'hb5)) ?
              wire1252 : wire1250[(5'h10):(4'hd)]))) ?
          reg1255[(4'hb):(4'ha)] : $signed(wire1250[(4'ha):(4'ha)]));
      for (forvar1259 = (1'h0); (forvar1259 < (1'h0)); forvar1259 = (forvar1259 + (1'h1)))
        begin
          reg1260 = $signed(forvar1259[(1'h1):(1'h1)]);
          reg1261 <= reg1256[(2'h2):(2'h2)];
        end
      reg1262 <= (~|$unsigned($signed(((reg1255 ? (7'h42) : wire1252) ?
          (reg1253 ? wire1252 : reg1254) : (&reg1261)))));
    end
  assign wire1263 = $signed($unsigned({reg1260[(4'he):(3'h6)], (!wire1257)}));
  assign wire1264 = (($unsigned(wire1251) > (($unsigned(reg1253) ?
                            (~^reg1255) : (7'h44)) && ((wire1257 < reg1262) ?
                            $unsigned(wire1263) : {wire1251}))) ?
                        $signed((($unsigned(wire1251) && $signed(reg1256)) + ({wire1257} ?
                            $signed(reg1262) : $unsigned((8'ha3))))) : (reg1260[(1'h0):(1'h0)] <<< (~|wire1257[(1'h1):(1'h0)])));
  always
    @(posedge clk) begin
      for (forvar1265 = (1'h0); (forvar1265 < (2'h2)); forvar1265 = (forvar1265 + (1'h1)))
        begin
          reg1266 = (wire1251[(1'h0):(1'h0)] ?
              $unsigned((($unsigned(reg1260) ?
                  $unsigned(forvar1259) : wire1264) <= (((8'hbe) && reg1255) ?
                  $unsigned(reg1253) : (wire1257 ?
                      reg1258 : (8'haa))))) : (8'haf));
          reg1267 <= wire1263;
          reg1268 = (+((8'hba) + wire1251[(4'hc):(4'hb)]));
          reg1269 <= (^~((8'haa) ?
              $signed(($unsigned(wire1249) >>> (reg1255 ?
                  reg1254 : wire1257))) : (reg1254 <<< (^wire1250))));
          reg1270 <= {$unsigned(reg1266[(3'h6):(2'h2)]),
              ((~&$signed(wire1251)) ?
                  ($unsigned(reg1266[(3'h6):(2'h2)]) ?
                      reg1261[(3'h6):(2'h3)] : $unsigned($unsigned(reg1260))) : reg1260)};
        end
    end
  always
    @(posedge clk) begin
      reg1271 <= ($unsigned((wire1252[(2'h2):(1'h1)] << ((reg1261 >>> (8'ha1)) <= (wire1250 ^~ reg1256)))) & (~^(-wire1251)));
    end
  assign wire1272 = wire1251;
  always
    @(posedge clk) begin
      reg1273 = ((((reg1266 <= reg1262) << $signed($signed((8'ha5)))) ?
          reg1269 : $unsigned((~|(reg1266 ?
              (8'ha8) : forvar1259)))) < (($signed((forvar1265 ?
          wire1252 : reg1266)) ^~ ((|wire1257) && $signed(wire1249))) << (8'hac)));
      reg1274 = (^~reg1269[(5'h10):(2'h2)]);
      reg1275 <= $signed({($unsigned(reg1254) - reg1268[(3'h7):(1'h1)]),
          $unsigned(wire1250)});
    end
  always
    @(posedge clk) begin
      for (forvar1276 = (1'h0); (forvar1276 < (1'h1)); forvar1276 = (forvar1276 + (1'h1)))
        begin
          for (forvar1277 = (1'h0); (forvar1277 < (1'h1)); forvar1277 = (forvar1277 + (1'h1)))
            begin
              reg1278 = (^~wire1252[(1'h1):(1'h0)]);
              reg1279 <= {(~|$unsigned($signed(((8'hbf) > reg1273)))),
                  (reg1267[(2'h3):(1'h1)] ?
                      {$signed((reg1260 && reg1270)),
                          reg1278[(2'h2):(1'h0)]} : ($signed($unsigned(reg1278)) ?
                          $signed($unsigned(reg1273)) : {$signed(reg1253),
                              reg1274}))};
              reg1280 <= (&{({wire1252} ?
                      forvar1265[(4'h9):(3'h6)] : $signed({reg1253})),
                  reg1271[(1'h0):(1'h0)]});
              reg1281 <= $signed($unsigned((^~(8'hbe))));
            end
          reg1282 <= ({$signed(forvar1276[(4'h8):(3'h6)])} - reg1274);
          reg1283 <= {(!(wire1257 | (reg1274[(1'h1):(1'h1)] + reg1268)))};
        end
      reg1284 <= $unsigned(forvar1276);
      reg1285 = ($unsigned(reg1274) ?
          $unsigned(reg1256[(4'h9):(3'h7)]) : (wire1252 ?
              {($unsigned((8'ha3)) * {reg1255, reg1256}),
                  reg1278[(3'h5):(1'h1)]} : $signed(((wire1251 ?
                      reg1283 : reg1271) ?
                  (wire1250 != reg1284) : forvar1265[(4'h8):(1'h0)]))));
    end
  assign wire1286 = (8'ha7);
  always
    @(posedge clk) begin
      reg1287 <= {(reg1271[(3'h7):(3'h7)] > $unsigned($unsigned(reg1256)))};
      for (forvar1288 = (1'h0); (forvar1288 < (2'h3)); forvar1288 = (forvar1288 + (1'h1)))
        begin
          reg1289 <= ((+$unsigned(($unsigned(wire1250) ?
              reg1271 : forvar1259[(1'h1):(1'h0)]))) <<< forvar1265);
        end
      reg1290 <= $signed(((reg1282[(4'ha):(4'h8)] ?
          {(forvar1259 ? forvar1288 : reg1273),
              $signed(reg1282)} : $unsigned({reg1285})) ^~ ($unsigned(reg1279[(2'h3):(1'h0)]) ?
          reg1270 : $unsigned($signed(reg1271)))));
    end
  assign wire1291 = $unsigned({(8'hb8),
                        (|{wire1264, wire1263[(5'h10):(2'h2)]})});
  always
    @(posedge clk) begin
      reg1292 <= (8'ha0);
    end
  always
    @(posedge clk) begin
      reg1293 <= ((^wire1249) ?
          wire1291 : $unsigned(({$signed(reg1285), reg1273[(1'h1):(1'h1)]} ?
              ((8'ha9) ?
                  wire1249[(4'h9):(3'h7)] : $unsigned(wire1251)) : $signed((wire1252 >>> reg1266)))));
      reg1294 <= $signed({wire1272,
          (~($signed(wire1272) && reg1258[(4'hf):(4'hd)]))});
      reg1295 = $unsigned(reg1285[(1'h1):(1'h0)]);
      reg1296 <= $unsigned({reg1261});
    end
  assign wire1297 = (^~((((reg1255 ?
                            reg1285 : forvar1288) > reg1254[(2'h3):(1'h1)]) ?
                        reg1267[(3'h7):(3'h4)] : {(reg1278 || reg1256)}) ^~ $unsigned({reg1281[(1'h1):(1'h0)],
                        $unsigned(reg1273)})));
  assign wire1298 = (reg1294 ?
                        $unsigned(forvar1276) : ({(8'hbe),
                            (8'haf)} + $unsigned(reg1296)));
  always
    @(posedge clk) begin
      reg1299 <= (reg1274[(1'h0):(1'h0)] != ({wire1291[(1'h0):(1'h0)],
          reg1290} <= ($signed($unsigned((8'ha0))) > ((reg1275 <= (8'ha5)) ^~ (^wire1249)))));
      reg1300 <= $signed($signed($unsigned((!$signed((8'ha2))))));
    end
  assign wire1301 = {$signed($unsigned(((!reg1283) ?
                            forvar1276[(2'h3):(2'h2)] : {wire1264, (8'hb9)}))),
                        $unsigned($signed(wire1291[(3'h4):(1'h0)]))};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1186
#( parameter param1240 = {(~|((~^((8'hb6) ? (8'hb0) : (8'hb0))) >> ((8'h9d) ? ((8'ha7) <= (8'h9e)) : {(7'h40)})))} )
(y, clk, wire1191, wire1190, wire1189, wire1188, wire1187);
  output wire [(32'h267):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire1191;
  input wire signed [(3'h6):(1'h0)] wire1190;
  input wire [(2'h2):(1'h0)] wire1189;
  input wire [(5'h15):(1'h0)] wire1188;
  input wire [(3'h4):(1'h0)] wire1187;
  reg signed [(4'hf):(1'h0)] reg1239 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1238 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1237 = (1'h0);
  reg [(3'h6):(1'h0)] reg1236 = (1'h0);
  reg [(4'hc):(1'h0)] reg1235 = (1'h0);
  reg [(4'hf):(1'h0)] reg1233 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1234 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1233 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1232 = (1'h0);
  reg [(4'h9):(1'h0)] reg1231 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1230 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1229 = (1'h0);
  reg [(4'h8):(1'h0)] reg1228 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1227 = (1'h0);
  reg [(2'h2):(1'h0)] reg1226 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1225 = (1'h0);
  reg [(4'h8):(1'h0)] reg1224 = (1'h0);
  reg [(4'he):(1'h0)] reg1223 = (1'h0);
  wire [(5'h13):(1'h0)] wire1222;
  reg [(5'h13):(1'h0)] reg1221 = (1'h0);
  reg [(4'hf):(1'h0)] reg1220 = (1'h0);
  reg [(4'hf):(1'h0)] reg1219 = (1'h0);
  reg [(5'h15):(1'h0)] reg1218 = (1'h0);
  reg [(3'h6):(1'h0)] reg1217 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1216 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1215 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1214 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1213 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1212 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1211 = (1'h0);
  reg [(5'h15):(1'h0)] reg1210 = (1'h0);
  reg [(4'he):(1'h0)] reg1209 = (1'h0);
  wire [(5'h14):(1'h0)] wire1208;
  wire signed [(5'h11):(1'h0)] wire1207;
  wire signed [(5'h14):(1'h0)] wire1206;
  reg [(4'hf):(1'h0)] reg1205 = (1'h0);
  reg [(5'h11):(1'h0)] reg1204 = (1'h0);
  wire [(4'hc):(1'h0)] wire1203;
  reg [(3'h6):(1'h0)] reg1202 = (1'h0);
  reg [(3'h6):(1'h0)] reg1201 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1200 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1199 = (1'h0);
  reg [(4'ha):(1'h0)] reg1198 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire1197;
  reg signed [(3'h6):(1'h0)] reg1196 = (1'h0);
  reg [(2'h3):(1'h0)] reg1195 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1194 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1193 = (1'h0);
  wire [(3'h5):(1'h0)] wire1192;
  assign y = {reg1239,
                 reg1238,
                 forvar1237,
                 reg1236,
                 reg1235,
                 reg1233,
                 reg1234,
                 forvar1233,
                 reg1232,
                 reg1231,
                 reg1230,
                 reg1229,
                 reg1228,
                 forvar1227,
                 reg1226,
                 reg1225,
                 reg1224,
                 reg1223,
                 wire1222,
                 reg1221,
                 reg1220,
                 reg1219,
                 reg1218,
                 reg1217,
                 reg1216,
                 forvar1215,
                 reg1214,
                 reg1213,
                 reg1212,
                 forvar1211,
                 reg1210,
                 reg1209,
                 wire1208,
                 wire1207,
                 wire1206,
                 reg1205,
                 reg1204,
                 wire1203,
                 reg1202,
                 reg1201,
                 reg1200,
                 reg1199,
                 reg1198,
                 wire1197,
                 reg1196,
                 reg1195,
                 forvar1194,
                 reg1193,
                 wire1192,
                 (1'h0)};
  assign wire1192 = $unsigned(($signed(wire1187) | (~wire1189)));
  always
    @(posedge clk) begin
      reg1193 = wire1189[(1'h0):(1'h0)];
      for (forvar1194 = (1'h0); (forvar1194 < (3'h4)); forvar1194 = (forvar1194 + (1'h1)))
        begin
          reg1195 <= (&((&$unsigned({wire1188,
              wire1188})) ~^ wire1190[(3'h6):(3'h4)]));
        end
      reg1196 = ({wire1189[(1'h1):(1'h0)],
              ($unsigned(forvar1194) ?
                  (reg1193[(3'h7):(2'h3)] ?
                      (forvar1194 ?
                          wire1192 : wire1192) : (!wire1192)) : (^~$unsigned(wire1191)))} ?
          ((8'hbc) ?
              ($unsigned(wire1192) ?
                  $unsigned($unsigned(reg1195)) : (~^wire1187[(2'h2):(1'h1)])) : ((wire1188[(4'ha):(2'h2)] ^ $unsigned(wire1190)) ?
                  $unsigned(forvar1194) : ($signed((8'hbb)) ?
                      (-wire1190) : (wire1189 - wire1189)))) : (|wire1187[(3'h4):(1'h0)]));
    end
  assign wire1197 = {$unsigned(wire1187)};
  always
    @(posedge clk) begin
      reg1198 <= ($signed(($unsigned(wire1188) << wire1189[(1'h0):(1'h0)])) ?
          (reg1196[(3'h6):(1'h1)] * (wire1197 ?
              {wire1197[(4'hc):(4'hb)],
                  wire1192[(1'h1):(1'h1)]} : ((wire1187 == wire1189) ^ (wire1189 << wire1191)))) : (&(|wire1188)));
    end
  always
    @(posedge clk) begin
      reg1199 <= $unsigned(((forvar1194[(3'h4):(3'h4)] + (^(forvar1194 ?
              reg1193 : reg1198))) ?
          $unsigned((((8'hb4) ?
              forvar1194 : reg1196) <= $signed((8'hba)))) : ((~|$signed(wire1190)) ?
              (+{(8'hb4), wire1187}) : reg1196)));
      reg1200 <= $unsigned((8'hb3));
      reg1201 <= (reg1193[(4'h8):(2'h3)] ?
          $unsigned(wire1187[(1'h1):(1'h0)]) : $signed((&wire1190[(3'h6):(3'h6)])));
      reg1202 <= reg1200[(2'h2):(2'h2)];
    end
  assign wire1203 = $unsigned((8'ha5));
  always
    @(posedge clk) begin
      reg1204 <= {$signed((((wire1191 ? reg1193 : reg1199) < $signed(reg1193)) ?
              ({wire1191, wire1187} | (8'hb0)) : reg1199)),
          $signed((reg1202 ?
              (&(wire1188 >>> wire1189)) : reg1199[(2'h3):(2'h3)]))};
      reg1205 <= forvar1194[(2'h2):(1'h0)];
    end
  assign wire1206 = (($signed((~$signed(reg1199))) || ($unsigned($signed((8'ha8))) > $signed(reg1195[(1'h1):(1'h1)]))) != $signed(reg1201));
  assign wire1207 = $unsigned(wire1206);
  assign wire1208 = $unsigned($signed({(wire1206[(4'hd):(4'h9)] ?
                            wire1203 : wire1206[(4'ha):(2'h2)]),
                        ($signed(reg1198) < {wire1189, (8'h9c)})}));
  always
    @(posedge clk) begin
      reg1209 <= wire1191[(5'h13):(3'h4)];
      reg1210 <= wire1192;
    end
  always
    @(posedge clk) begin
      for (forvar1211 = (1'h0); (forvar1211 < (2'h2)); forvar1211 = (forvar1211 + (1'h1)))
        begin
          reg1212 = ((~reg1198) ?
              (reg1204 << (^~reg1200[(1'h0):(1'h0)])) : ((reg1198 << {(^reg1200),
                  $unsigned(reg1195)}) >>> reg1209[(1'h1):(1'h0)]));
          reg1213 <= (|(!(|$signed(reg1198))));
          reg1214 <= $unsigned(reg1213);
          for (forvar1215 = (1'h0); (forvar1215 < (1'h1)); forvar1215 = (forvar1215 + (1'h1)))
            begin
              reg1216 <= $unsigned(reg1198);
              reg1217 <= (-$signed(reg1214[(4'h9):(3'h7)]));
              reg1218 <= $unsigned((~((((8'hab) - wire1207) ^~ (reg1217 ^~ reg1201)) ?
                  wire1203[(3'h4):(2'h3)] : ($signed((7'h44)) ?
                      (forvar1211 ? reg1202 : (8'haa)) : wire1188))));
              reg1219 <= (reg1212[(1'h1):(1'h0)] ?
                  {({$unsigned(reg1202)} ?
                          reg1196[(3'h6):(3'h5)] : (wire1207[(3'h5):(3'h5)] != {reg1201,
                              forvar1215}))} : $signed(($signed($signed(wire1203)) ?
                      {(wire1188 ?
                              wire1208 : (8'hbb))} : (^~$signed(reg1205)))));
              reg1220 = $signed(forvar1194);
            end
          reg1221 = $unsigned(wire1203[(4'ha):(4'h8)]);
        end
    end
  assign wire1222 = wire1208[(2'h2):(2'h2)];
  always
    @(posedge clk) begin
      reg1223 <= (-reg1214[(3'h4):(2'h3)]);
      reg1224 <= (~|(reg1202[(1'h0):(1'h0)] <= (~(&(7'h41)))));
      reg1225 = $unsigned($signed(($signed((wire1191 | wire1190)) + $unsigned(wire1187[(3'h4):(1'h1)]))));
      reg1226 <= $signed({(((8'ha0) ? (|(7'h42)) : reg1218[(4'ha):(3'h6)]) ?
              {(~&reg1212)} : (reg1221 << ((7'h42) ? forvar1211 : reg1204))),
          ({(|reg1210), {reg1220}} >= forvar1194)});
    end
  always
    @(posedge clk) begin
      for (forvar1227 = (1'h0); (forvar1227 < (3'h4)); forvar1227 = (forvar1227 + (1'h1)))
        begin
          reg1228 <= $signed($unsigned(wire1222[(5'h13):(4'h8)]));
          reg1229 = (wire1203 ?
              ((reg1199[(4'h8):(1'h0)] ?
                  ($unsigned(reg1224) ?
                      $signed(wire1191) : wire1188) : ((&wire1222) ?
                      (reg1204 == (8'hb9)) : (reg1220 & wire1188))) == wire1206) : ((|{reg1193}) ?
                  $unsigned((((8'ha8) ? reg1204 : reg1220) ?
                      (forvar1194 == reg1198) : wire1208[(3'h4):(1'h0)])) : ({reg1223[(3'h4):(2'h2)],
                      (reg1228 ? forvar1215 : forvar1215)} >> (^(~|reg1216)))));
          reg1230 <= wire1206;
          reg1231 <= reg1225;
          reg1232 <= reg1220[(1'h1):(1'h1)];
        end
      if (reg1231)
        begin
          for (forvar1233 = (1'h0); (forvar1233 < (3'h4)); forvar1233 = (forvar1233 + (1'h1)))
            begin
              reg1234 <= ($unsigned(({reg1212} ?
                  $unsigned(reg1228) : wire1192)) - (-reg1196));
            end
        end
      else
        begin
          reg1233 = {($signed(wire1208[(3'h5):(2'h3)]) - (reg1202 ?
                  $unsigned($unsigned(reg1220)) : reg1193))};
          reg1234 <= ((~|$signed((reg1221[(2'h2):(1'h1)] != $unsigned(reg1223)))) ?
              {$unsigned($signed(reg1232))} : (((~&reg1225) + reg1234) ?
                  $unsigned(reg1216[(3'h7):(1'h1)]) : (((-wire1189) && (reg1221 ?
                          reg1219 : reg1216)) ?
                      wire1188 : ($signed((8'ha3)) * $unsigned(reg1199)))));
          reg1235 <= {(reg1205 ?
                  (($signed(reg1209) ?
                      wire1191[(4'h9):(4'h9)] : $signed(forvar1227)) <<< (~&(!reg1218))) : $unsigned((^(reg1198 ?
                      reg1193 : (8'ha5))))),
              (~|(((!forvar1233) ?
                  (-wire1189) : $unsigned(wire1208)) - reg1232))};
        end
      reg1236 <= reg1201;
      for (forvar1237 = (1'h0); (forvar1237 < (2'h2)); forvar1237 = (forvar1237 + (1'h1)))
        begin
          reg1238 <= ((&reg1217[(2'h2):(1'h1)]) ?
              $signed(forvar1227) : $unsigned((&$signed($unsigned(reg1199)))));
        end
      reg1239 <= $unsigned((wire1222 > (-$unsigned(reg1216))));
    end
endmodule