(* use_dsp48="no" *) (* use_dsp="no" *) module top
#( parameter param210 = (~&(~|(({(8'ha4), (7'h42)} - ((8'ha5) <<< (8'hb9))) < (((8'h9f) < (8'h9e)) ? (8'hbf) : (|(8'ha9))))))
, parameter param211 = param210 )
(y, clk, wire0, wire1, wire2, wire3);
  output wire [(32'h2b6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h3):(1'h0)] wire0;
  input wire [(4'hc):(1'h0)] wire1;
  input wire signed [(2'h3):(1'h0)] wire2;
  input wire signed [(4'hb):(1'h0)] wire3;
  reg signed [(4'hd):(1'h0)] reg209 = (1'h0);
  reg [(5'h13):(1'h0)] reg208 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg207 = (1'h0);
  wire [(4'h9):(1'h0)] wire198;
  wire [(5'h13):(1'h0)] wire197;
  wire [(5'h15):(1'h0)] wire196;
  wire [(4'hc):(1'h0)] wire195;
  reg [(4'hb):(1'h0)] reg4 = (1'h0);
  wire [(4'h8):(1'h0)] wire5;
  wire signed [(4'hf):(1'h0)] wire6;
  reg signed [(4'ha):(1'h0)] reg7 = (1'h0);
  reg [(4'ha):(1'h0)] reg8 = (1'h0);
  reg [(5'h13):(1'h0)] reg9 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg10 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg11 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg12 = (1'h0);
  reg [(2'h2):(1'h0)] reg13 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg14 = (1'h0);
  reg [(5'h13):(1'h0)] reg15 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg16 = (1'h0);
  reg [(5'h13):(1'h0)] reg17 = (1'h0);
  reg [(4'hc):(1'h0)] reg18 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg19 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg20 = (1'h0);
  reg [(2'h3):(1'h0)] reg21 = (1'h0);
  reg [(5'h13):(1'h0)] reg22 = (1'h0);
  reg [(4'ha):(1'h0)] reg23 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg24 = (1'h0);
  reg [(5'h15):(1'h0)] reg25 = (1'h0);
  reg [(4'h9):(1'h0)] reg26 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg27 = (1'h0);
  reg [(3'h7):(1'h0)] reg28 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg29 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg30 = (1'h0);
  reg [(5'h11):(1'h0)] reg31 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg32 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg33 = (1'h0);
  reg [(5'h15):(1'h0)] reg34 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg35 = (1'h0);
  reg [(5'h15):(1'h0)] reg36 = (1'h0);
  reg [(5'h10):(1'h0)] reg37 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg38 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire39;
  wire [(5'h14):(1'h0)] wire155;
  wire [(4'hd):(1'h0)] wire157;
  wire [(4'hd):(1'h0)] wire158;
  wire signed [(4'hc):(1'h0)] wire193;
  wire [(4'h8):(1'h0)] wire200;
  wire [(3'h4):(1'h0)] wire201;
  wire signed [(3'h6):(1'h0)] wire202;
  wire [(5'h11):(1'h0)] wire203;
  wire signed [(4'h8):(1'h0)] wire205;
  assign y = {reg209,
                 reg208,
                 reg207,
                 wire198,
                 wire197,
                 wire196,
                 wire195,
                 reg4,
                 wire5,
                 wire6,
                 reg7,
                 reg8,
                 reg9,
                 reg10,
                 reg11,
                 reg12,
                 reg13,
                 reg14,
                 reg15,
                 reg16,
                 reg17,
                 reg18,
                 reg19,
                 reg20,
                 reg21,
                 reg22,
                 reg23,
                 reg24,
                 reg25,
                 reg26,
                 reg27,
                 reg28,
                 reg29,
                 reg30,
                 reg31,
                 reg32,
                 reg33,
                 reg34,
                 reg35,
                 reg36,
                 reg37,
                 reg38,
                 wire39,
                 wire155,
                 wire157,
                 wire158,
                 wire193,
                 wire200,
                 wire201,
                 wire202,
                 wire203,
                 wire205,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg4 <= (^~(~(-$signed($unsigned((8'hab))))));
    end
  assign wire5 = (&{{(reg4[(2'h3):(1'h0)] >> $unsigned(reg4)),
                         ((wire0 == wire2) ~^ wire3)}});
  assign wire6 = wire5;
  always
    @(posedge clk) begin
      reg7 <= {($signed((8'hb1)) ?
              ((8'ha0) & wire6[(1'h0):(1'h0)]) : ((reg4[(3'h7):(3'h6)] ?
                      ((8'ha0) ? wire5 : reg4) : (wire0 + reg4)) ?
                  wire3 : $unsigned($unsigned(wire1))))};
      reg8 <= $signed(wire6[(4'hf):(1'h0)]);
      reg9 <= $unsigned($signed(wire2));
      reg10 <= wire6[(1'h1):(1'h0)];
      reg11 <= $unsigned(reg4[(2'h3):(1'h1)]);
    end
  always
    @(posedge clk) begin
      if ($unsigned(reg9[(1'h1):(1'h1)]))
        begin
          reg12 <= reg11;
        end
      else
        begin
          if (wire5[(1'h0):(1'h0)])
            begin
              reg12 <= $unsigned($unsigned(($unsigned(reg10) + ({(8'ha2),
                  reg10} * $unsigned(reg4)))));
              reg13 <= wire5[(2'h3):(2'h2)];
            end
          else
            begin
              reg12 <= ($unsigned($signed($unsigned((7'h44)))) ?
                  (~^$unsigned($signed((reg13 | (8'ha9))))) : {$unsigned(($signed(reg8) * wire5[(2'h3):(1'h1)]))});
              reg13 <= $signed({{wire6[(4'he):(1'h0)]}, reg8});
              reg14 <= reg13;
            end
          reg15 <= wire0;
          reg16 <= reg11[(1'h1):(1'h0)];
          reg17 <= ((^(^$signed((~wire0)))) ?
              {reg8[(4'ha):(2'h3)],
                  $signed((reg10 ?
                      reg11[(1'h0):(1'h0)] : {reg8,
                          wire3}))} : (((~|reg7) << (+(8'ha1))) ?
                  wire2[(2'h3):(1'h1)] : reg13[(2'h2):(2'h2)]));
        end
      if ({$signed(wire6), $unsigned(reg13[(1'h0):(1'h0)])})
        begin
          if (((+({reg17} || (~^(wire2 ? reg11 : wire5)))) ?
              ((((8'hbe) ^~ wire5[(2'h2):(2'h2)]) * reg10[(3'h5):(1'h1)]) ^ reg10) : $unsigned((&((~reg10) + wire0)))))
            begin
              reg18 <= {reg14};
              reg19 <= (+wire5[(1'h0):(1'h0)]);
              reg20 <= (~$signed(($unsigned((&reg17)) ^ (8'ha2))));
              reg21 <= (~((((wire1 ? reg4 : reg20) ? $signed(reg8) : reg15) ?
                  {(~reg18), $unsigned(reg7)} : (wire0 ?
                      reg12 : reg9)) != {$unsigned((reg14 ? reg14 : (8'haf))),
                  $signed((+wire2))}));
            end
          else
            begin
              reg18 <= $signed($unsigned((reg19[(3'h6):(1'h1)] ?
                  reg10[(3'h6):(1'h0)] : reg11[(2'h2):(1'h1)])));
              reg19 <= (reg20[(3'h7):(3'h5)] >= reg21);
              reg20 <= $signed((reg20[(2'h3):(2'h3)] ?
                  reg20[(1'h0):(1'h0)] : ($signed((reg20 << reg8)) ?
                      wire6[(3'h4):(2'h3)] : $unsigned((reg14 ?
                          reg12 : wire2)))));
              reg21 <= $unsigned((reg17 && $signed((reg17[(4'hd):(3'h4)] <= $signed((8'ha5))))));
              reg22 <= (|reg8);
            end
          if (wire3)
            begin
              reg23 <= {wire5};
              reg24 <= $unsigned((reg10 && (($signed(reg10) ?
                  $unsigned(reg11) : wire0) <<< reg20[(4'h9):(3'h5)])));
            end
          else
            begin
              reg23 <= (reg7 + (reg16[(3'h7):(3'h7)] <<< {reg11, reg23}));
              reg24 <= ((($signed($signed((8'hb0))) <= $unsigned((wire5 | wire5))) ?
                  {reg12[(4'hc):(4'hc)]} : reg12) <= wire0);
              reg25 <= $unsigned($signed({(+{reg10, reg11}),
                  (wire3[(3'h6):(2'h3)] ?
                      $signed(reg21) : ((8'hb6) ? reg18 : reg21))}));
              reg26 <= reg15[(3'h5):(1'h1)];
            end
          reg27 <= ($signed(wire3[(1'h1):(1'h1)]) ?
              reg12 : (($unsigned((reg11 | wire6)) >>> (reg14[(3'h7):(1'h1)] ?
                  (wire1 ? wire3 : reg17) : $unsigned(reg18))) && reg22));
        end
      else
        begin
          reg18 <= ((+$signed($unsigned((^reg22)))) ?
              $signed(wire1) : ($unsigned(reg20) ?
                  (($unsigned(reg23) + reg7) | ((reg21 <<< reg14) > reg27[(3'h6):(3'h6)])) : $unsigned($signed($signed((8'hb0))))));
          if (($signed(wire0) ?
              $unsigned($unsigned($unsigned($signed(reg25)))) : $unsigned(reg18[(3'h6):(3'h4)])))
            begin
              reg19 <= reg8[(3'h4):(2'h3)];
              reg20 <= reg27;
            end
          else
            begin
              reg19 <= $unsigned($unsigned(reg10[(4'h8):(3'h4)]));
              reg20 <= $signed(($signed(reg20[(3'h5):(2'h3)]) >= reg24));
              reg21 <= ((($signed($unsigned(wire0)) ^ $unsigned((reg13 ?
                      wire3 : wire5))) ?
                  (reg8 <<< (reg20[(1'h1):(1'h0)] >> wire3[(1'h1):(1'h1)])) : ($unsigned(wire0[(2'h3):(1'h1)]) ?
                      ((reg8 > (8'hba)) >>> (+reg8)) : (~&{reg14,
                          (8'hba)}))) >> (reg9[(1'h1):(1'h1)] + wire2));
              reg22 <= (~$signed(reg25));
            end
          reg23 <= (8'ha9);
          reg24 <= ($signed(reg7[(2'h3):(1'h0)]) ?
              $signed($unsigned(((wire1 != (8'hb2)) ?
                  (reg27 ? reg8 : reg14) : (reg23 & reg24)))) : (({(reg24 ?
                          wire5 : reg22)} ?
                  $unsigned(wire2[(1'h0):(1'h0)]) : $unsigned(reg26)) ^ wire1));
          reg25 <= (({reg12} ?
              ((-wire5) != ($unsigned(reg12) ?
                  (reg20 ~^ reg21) : (reg8 <= reg8))) : {reg23[(1'h0):(1'h0)],
                  reg18}) >= (wire6 ?
              $signed(($signed(wire2) ?
                  (wire5 * reg23) : reg15)) : ($signed({reg26}) & $unsigned((~^reg15)))));
        end
      reg28 <= (^~reg14);
      if ({$unsigned($unsigned(reg8))})
        begin
          reg29 <= wire2;
        end
      else
        begin
          if ($signed((reg10[(2'h3):(2'h2)] | reg4)))
            begin
              reg29 <= $unsigned($unsigned($signed((~(reg13 ?
                  reg11 : reg20)))));
              reg30 <= ((!(^(^~wire2))) ?
                  ({{(~^wire1)},
                      $signed($signed((8'hbe)))} ^ $signed((8'hb4))) : reg4);
              reg31 <= reg22;
              reg32 <= {($unsigned((^~(reg16 <<< wire2))) ?
                      (+reg14) : (-$unsigned(reg14)))};
              reg33 <= ($signed(reg10[(4'h9):(3'h6)]) ?
                  reg11[(3'h5):(3'h5)] : $unsigned(reg9[(2'h2):(2'h2)]));
            end
          else
            begin
              reg29 <= reg14;
              reg30 <= $unsigned(reg14);
              reg31 <= reg31;
              reg32 <= (8'hbe);
              reg33 <= (reg4[(3'h4):(2'h3)] ?
                  reg14 : (((((8'hbf) ? reg26 : wire6) ?
                          (8'haf) : (~&reg33)) ~^ ({(7'h40),
                          reg31} - (^~reg11))) ?
                      $signed((~&$unsigned((8'hbb)))) : reg25[(3'h4):(3'h4)]));
            end
          reg34 <= $unsigned(reg19);
          if ({(reg32 ?
                  (reg24[(4'he):(3'h4)] ?
                      ((!reg34) ?
                          (&(8'h9c)) : {reg18}) : $signed($unsigned((8'ha5)))) : {reg20[(1'h0):(1'h0)],
                      reg23[(3'h4):(1'h0)]}),
              ({wire1[(3'h6):(1'h1)]} ? reg23 : {reg22[(3'h5):(1'h1)]})})
            begin
              reg35 <= (|$unsigned($signed(((-wire2) > reg26))));
              reg36 <= reg12[(4'h8):(3'h4)];
              reg37 <= (((wire6 - reg33) ?
                      $signed($signed($unsigned(reg33))) : $unsigned($unsigned($signed(reg34)))) ?
                  ((8'hbb) ?
                      (8'ha8) : reg36[(3'h5):(1'h1)]) : ((-$unsigned((reg23 ?
                      reg36 : reg24))) >> $signed((|$unsigned((8'hab))))));
              reg38 <= reg22;
            end
          else
            begin
              reg35 <= (^$unsigned(($unsigned(reg19) | $unsigned(wire0[(2'h3):(1'h0)]))));
              reg36 <= reg35[(4'ha):(4'h8)];
              reg37 <= $unsigned(reg10[(4'h9):(1'h0)]);
            end
        end
    end
  assign wire39 = (~^(((^~(|(8'ha4))) ^~ {(+reg10)}) ?
                      $signed(({reg8, (8'ha4)} | (reg30 ?
                          reg29 : reg33))) : reg25));
  module40 modinst156 (.wire42(reg24), .wire44(reg9), .wire43(wire1), .wire41(reg18), .clk(clk), .y(wire155));
  assign wire157 = (|$unsigned((~&((8'hac) >= (wire1 ? reg32 : reg15)))));
  assign wire158 = $signed(({(^~(reg27 ?
                           reg4 : reg28))} <<< $signed((~|{(8'hb5)}))));
  module159 modinst194 (.y(wire193), .clk(clk), .wire161(reg19), .wire164(reg30), .wire160(reg37), .wire162(reg10), .wire163(reg36));
  assign wire195 = {((8'hb9) * $unsigned(reg16)), reg22[(5'h12):(2'h2)]};
  assign wire196 = (wire6 ?
                       {(reg17 ?
                               (8'hb2) : $unsigned(reg35))} : $unsigned({(8'hbf),
                           {(reg20 >= wire2), $signed(wire3)}}));
  assign wire197 = (wire3 ?
                       wire1 : $unsigned((|((reg27 ? reg32 : wire5) ?
                           (reg4 ^ reg9) : (reg37 <<< (8'haf))))));
  module46 modinst199 (.wire50(reg23), .wire51(reg4), .wire48(reg14), .y(wire198), .wire47(reg7), .wire49(reg31), .clk(clk));
  assign wire200 = $unsigned($signed({(~^$unsigned((8'hba))),
                       $unsigned((|(8'h9e)))}));
  assign wire201 = (^~(^(^((reg4 | (8'h9f)) ?
                       (reg8 - (7'h41)) : (reg33 ? (7'h44) : wire155)))));
  assign wire202 = ($unsigned((|(reg32[(1'h0):(1'h0)] ?
                       $unsigned(wire5) : $signed(wire157)))) && wire39);
  module113 modinst204 (.wire115(reg26), .y(wire203), .wire117(reg30), .wire114(reg9), .clk(clk), .wire116(wire39));
  module88 modinst206 (.wire89(reg17), .wire90(reg28), .wire91(wire155), .y(wire205), .wire93(reg25), .clk(clk), .wire92(reg14));
  always
    @(posedge clk) begin
      reg207 <= (~^$signed(wire0));
      reg208 <= ($unsigned((|reg30[(3'h6):(3'h6)])) ?
          (|({$signed(reg37)} == $signed((&reg22)))) : wire205[(3'h6):(3'h5)]);
      reg209 <= ((wire6[(1'h0):(1'h0)] ?
              (~|$unsigned(((8'hbf) ?
                  wire1 : reg26))) : (reg208 >>> ($unsigned(reg35) ~^ $unsigned(wire6)))) ?
          reg21[(2'h2):(1'h1)] : ($signed(reg14[(5'h10):(4'he)]) < (((reg13 ?
                  reg14 : reg37) || $signed(wire3)) ?
              ((reg20 ? (8'ha4) : reg25) ?
                  $unsigned(wire198) : (reg7 ?
                      wire3 : reg23)) : (~(reg11 == reg23)))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module159
#( parameter param191 = ((!{(((7'h42) ? (8'ha3) : (8'h9c)) ? ((8'h9f) >>> (7'h44)) : (~|(8'ha1)))}) != ((^~(8'h9f)) ? ((|((7'h44) ? (8'hba) : (8'hb5))) <= (((8'ha0) ? (8'hb2) : (8'hb0)) ? ((8'hb1) ? (8'hbc) : (8'hba)) : ((8'ha7) ? (8'ha3) : (8'hae)))) : ({(!(8'had))} >> (~((8'ha4) >= (8'hab))))))
, parameter param192 = {(|(8'hae))} )
(y, clk, wire164, wire163, wire162, wire161, wire160);
  output wire [(32'h159):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire164;
  input wire signed [(5'h15):(1'h0)] wire163;
  input wire signed [(4'hc):(1'h0)] wire162;
  input wire [(4'h8):(1'h0)] wire161;
  input wire [(3'h6):(1'h0)] wire160;
  wire [(3'h5):(1'h0)] wire190;
  wire [(5'h12):(1'h0)] wire189;
  reg signed [(5'h12):(1'h0)] reg188 = (1'h0);
  reg [(2'h3):(1'h0)] reg187 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg186 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg185 = (1'h0);
  reg [(4'hf):(1'h0)] reg184 = (1'h0);
  reg [(4'h8):(1'h0)] reg183 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg182 = (1'h0);
  reg [(3'h5):(1'h0)] reg181 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg180 = (1'h0);
  reg [(4'h8):(1'h0)] reg179 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg178 = (1'h0);
  reg [(5'h14):(1'h0)] reg177 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg176 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg175 = (1'h0);
  reg [(5'h12):(1'h0)] reg174 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg173 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg172 = (1'h0);
  reg [(4'he):(1'h0)] reg171 = (1'h0);
  reg [(5'h10):(1'h0)] reg170 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire169;
  wire signed [(5'h15):(1'h0)] wire168;
  wire signed [(5'h15):(1'h0)] wire167;
  wire [(5'h13):(1'h0)] wire166;
  wire [(5'h12):(1'h0)] wire165;
  assign y = {wire190,
                 wire189,
                 reg188,
                 reg187,
                 reg186,
                 reg185,
                 reg184,
                 reg183,
                 reg182,
                 reg181,
                 reg180,
                 reg179,
                 reg178,
                 reg177,
                 reg176,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 reg171,
                 reg170,
                 wire169,
                 wire168,
                 wire167,
                 wire166,
                 wire165,
                 (1'h0)};
  assign wire165 = wire160[(3'h6):(3'h6)];
  assign wire166 = ($unsigned({$signed(((8'hb2) ?
                           wire165 : wire161))}) ^~ (+wire162));
  assign wire167 = ({wire166} ?
                       (~&wire166) : $signed((wire160[(1'h1):(1'h1)] ?
                           $unsigned(wire166) : $signed(wire166))));
  assign wire168 = wire167;
  assign wire169 = {wire161[(4'h8):(3'h4)]};
  always
    @(posedge clk) begin
      reg170 <= ({{{$signed(wire167), (wire160 ? wire163 : wire168)}},
              {{(~&wire164), (wire160 ? wire167 : wire165)}, wire161}} ?
          (~|(^$unsigned(((8'h9d) ? wire164 : wire166)))) : {(~&(&(wire169 ?
                  wire162 : wire160))),
              ($signed($unsigned((7'h43))) < (~&(wire161 ?
                  (8'haf) : (8'hbc))))});
      reg171 <= ({$unsigned({(~|wire163)}),
          ($signed((+wire161)) ^~ wire165)} <<< wire165[(4'hb):(4'h9)]);
      if ((((8'hb3) | (^wire165[(2'h3):(1'h1)])) ?
          $unsigned($unsigned(((wire161 < wire163) ?
              reg170[(3'h4):(2'h3)] : wire163))) : wire167))
        begin
          reg172 <= ((+((+$unsigned(wire162)) + ((wire161 ? wire166 : wire162) ?
              (~wire164) : $unsigned(wire163)))) ~^ ($signed($signed($unsigned((8'hab)))) ?
              (^(8'hb8)) : $signed((~|$unsigned(wire167)))));
          reg173 <= wire167;
          if (((~&wire161) ?
              (~(((|wire160) + wire160) >>> ($signed(wire163) ?
                  (reg173 ?
                      wire166 : wire164) : $signed((8'ha0))))) : $unsigned($unsigned({(wire162 ?
                      wire168 : wire165),
                  ((8'hbf) << reg170)}))))
            begin
              reg174 <= $signed($signed(wire168[(5'h10):(4'ha)]));
            end
          else
            begin
              reg174 <= $unsigned($signed($unsigned(wire169[(1'h1):(1'h1)])));
              reg175 <= ((($signed({wire163, wire160}) ?
                  $signed($unsigned(wire165)) : $unsigned((~(8'ha0)))) <= ($unsigned($signed(reg174)) >= $signed($signed(wire161)))) <<< wire160[(3'h4):(2'h3)]);
            end
          reg176 <= (((!$signed((wire169 * wire166))) ?
                  reg173 : (-$signed($signed(wire163)))) ?
              $signed(({wire164,
                  (&wire162)} ^ reg175)) : wire165[(4'he):(3'h7)]);
          reg177 <= $signed((wire164[(3'h4):(3'h4)] ?
              (|wire162) : reg174[(4'hd):(4'hc)]));
        end
      else
        begin
          reg172 <= wire168[(4'hd):(3'h4)];
          reg173 <= reg173;
          reg174 <= $signed((({{wire169,
                  wire162}} || (-reg171[(4'he):(4'ha)])) < (((~^reg176) && (reg177 < wire162)) ?
              $signed((wire161 ?
                  reg171 : reg177)) : (reg171 <<< (^~(8'h9d))))));
        end
      if ($signed(reg173))
        begin
          reg178 <= $unsigned((|{$signed($signed(wire167)),
              $unsigned((wire165 == reg170))}));
          if ($signed($signed(reg171)))
            begin
              reg179 <= $unsigned($signed((^reg174[(4'hb):(4'h8)])));
              reg180 <= (~(8'h9e));
            end
          else
            begin
              reg179 <= (reg175 ? wire166 : (!wire161[(3'h6):(2'h3)]));
              reg180 <= ((!$unsigned((!(wire165 ?
                  wire164 : wire169)))) < $unsigned(reg170[(2'h3):(2'h2)]));
              reg181 <= $unsigned(({(reg176 ?
                          $unsigned((8'ha9)) : (wire164 ? wire168 : (8'ha1)))} ?
                  $unsigned($unsigned($unsigned(reg174))) : (^~(reg171 ?
                      (~reg179) : (wire161 ? reg179 : reg179)))));
              reg182 <= (reg171[(4'ha):(2'h2)] == reg172);
            end
          reg183 <= (^(!$unsigned((7'h40))));
          if (reg175[(3'h4):(2'h2)])
            begin
              reg184 <= (^$signed(wire166[(4'he):(4'h8)]));
            end
          else
            begin
              reg184 <= (!$unsigned((({wire164, reg173} ?
                  $unsigned((8'hb2)) : reg181) * reg176[(3'h6):(3'h5)])));
              reg185 <= (-{wire169[(2'h2):(1'h0)]});
              reg186 <= ((~|({$signed(reg176)} ? wire168 : wire165)) ?
                  $signed($signed(((reg170 ?
                      wire167 : reg176) ^ (-reg171)))) : reg175);
            end
          if ($signed($signed(wire169)))
            begin
              reg187 <= (reg170[(4'h9):(3'h5)] ?
                  $unsigned((+$signed($unsigned(reg171)))) : (^((-(-reg184)) ^ (!reg176[(1'h0):(1'h0)]))));
            end
          else
            begin
              reg187 <= reg175;
            end
        end
      else
        begin
          reg178 <= {$signed(wire167[(4'hd):(2'h2)]),
              (reg170[(4'hd):(4'hc)] <<< $unsigned(wire165))};
          reg179 <= (reg184 ? $unsigned(reg177[(4'ha):(1'h0)]) : wire168);
          if (wire164)
            begin
              reg180 <= wire164[(4'ha):(3'h5)];
              reg181 <= ($signed($unsigned({$unsigned(reg185),
                  $unsigned(reg171)})) ~^ ($signed(reg171) ?
                  reg171[(4'h9):(4'h9)] : (&(8'hb1))));
            end
          else
            begin
              reg180 <= $signed(wire163[(3'h7):(3'h6)]);
              reg181 <= {$unsigned($signed(reg179)), wire164};
            end
          reg182 <= {$signed((~|(8'hbd))), $unsigned(wire166[(4'ha):(3'h5)])};
        end
      reg188 <= (reg179 ?
          (+((((8'hbd) < reg182) ?
              $unsigned((8'haa)) : wire165[(1'h1):(1'h1)]) << ($unsigned(reg187) ~^ reg182))) : wire169);
    end
  assign wire189 = ($signed(($unsigned((8'hae)) ~^ $signed((|wire163)))) * $unsigned(($unsigned((reg175 >> reg180)) ?
                       (reg172 ?
                           (wire167 ?
                               (8'haa) : reg186) : (-wire160)) : $signed($signed(reg188)))));
  assign wire190 = reg183[(3'h6):(3'h6)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module40
#( parameter param154 = (((8'hb4) ? ({(~&(8'ha0)), (&(8'h9d))} ? (((8'ha4) ? (8'hae) : (8'hb4)) ~^ {(8'ha5), (8'ha9)}) : (((8'had) < (8'hb9)) != ((8'hae) >> (8'hab)))) : {(8'ha6)}) <= (({((8'haf) & (8'ha1))} ? (-{(8'ha6), (8'ha5)}) : {(^(8'hb4)), ((8'hae) >>> (8'ha3))}) ? ((((8'ha7) > (8'hb0)) ? ((8'hbe) ? (8'ha3) : (8'haf)) : ((7'h43) & (8'ha6))) <<< (((8'had) * (7'h41)) ? ((8'haa) ^ (8'hb5)) : (|(8'hb3)))) : (((&(8'hbe)) || ((8'h9c) | (8'hb2))) ? {(&(8'h9c))} : (((8'ha9) ? (8'hba) : (8'hbe)) ^ (8'hbd))))) )
(y, clk, wire44, wire43, wire42, wire41);
  output wire [(32'h137):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire44;
  input wire signed [(4'hc):(1'h0)] wire43;
  input wire signed [(5'h14):(1'h0)] wire42;
  input wire [(4'hc):(1'h0)] wire41;
  wire signed [(4'hf):(1'h0)] wire153;
  wire [(4'hd):(1'h0)] wire152;
  wire signed [(3'h4):(1'h0)] wire151;
  wire [(3'h5):(1'h0)] wire150;
  wire signed [(3'h6):(1'h0)] wire149;
  reg signed [(4'hd):(1'h0)] reg148 = (1'h0);
  reg [(5'h10):(1'h0)] reg147 = (1'h0);
  reg [(4'h8):(1'h0)] reg146 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg145 = (1'h0);
  reg [(3'h5):(1'h0)] reg144 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg143 = (1'h0);
  reg signed [(4'he):(1'h0)] reg142 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg141 = (1'h0);
  reg [(3'h7):(1'h0)] reg140 = (1'h0);
  reg [(3'h4):(1'h0)] reg139 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg138 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire137;
  wire [(4'hc):(1'h0)] wire136;
  wire [(3'h4):(1'h0)] wire135;
  wire [(4'he):(1'h0)] wire134;
  wire signed [(5'h15):(1'h0)] wire133;
  wire [(3'h7):(1'h0)] wire131;
  wire signed [(2'h2):(1'h0)] wire112;
  wire [(4'hf):(1'h0)] wire111;
  wire signed [(3'h7):(1'h0)] wire110;
  wire [(4'h9):(1'h0)] wire109;
  wire [(4'h9):(1'h0)] wire108;
  wire [(5'h10):(1'h0)] wire86;
  wire signed [(5'h15):(1'h0)] wire45;
  wire [(3'h7):(1'h0)] wire106;
  assign y = {wire153,
                 wire152,
                 wire151,
                 wire150,
                 wire149,
                 reg148,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 reg143,
                 reg142,
                 reg141,
                 reg140,
                 reg139,
                 reg138,
                 wire137,
                 wire136,
                 wire135,
                 wire134,
                 wire133,
                 wire131,
                 wire112,
                 wire111,
                 wire110,
                 wire109,
                 wire108,
                 wire86,
                 wire45,
                 wire106,
                 (1'h0)};
  assign wire45 = {$signed(($signed(wire41[(3'h5):(3'h5)]) ^~ ((wire44 ?
                              wire41 : (8'hbd)) ?
                          (wire42 ? wire43 : (8'hb1)) : (-wire42)))),
                      $signed(wire44)};
  module46 modinst87 (wire86, clk, wire45, wire41, wire43, wire42, wire44);
  module88 modinst107 (wire106, clk, wire45, wire86, wire41, wire44, wire43);
  assign wire108 = wire106;
  assign wire109 = {{$signed(wire43[(4'h8):(1'h0)]),
                           $signed((((8'had) ^~ wire106) ?
                               (|wire42) : (wire43 ~^ wire41)))},
                       $signed(({wire106} ?
                           $unsigned((wire43 ?
                               wire108 : wire41)) : ($signed(wire108) ?
                               wire41[(3'h4):(1'h0)] : $unsigned(wire44))))};
  assign wire110 = ($unsigned($unsigned(((wire109 >>> wire44) > wire41[(4'h9):(4'h9)]))) ?
                       (^(&$signed(wire108))) : wire45);
  assign wire111 = (|(|(wire86 ?
                       $unsigned((8'hb5)) : $signed(wire106[(2'h3):(2'h2)]))));
  assign wire112 = ($unsigned(wire45) ? wire41 : wire43);
  module113 modinst132 (.clk(clk), .wire116(wire43), .wire114(wire44), .wire115(wire110), .y(wire131), .wire117(wire108));
  assign wire133 = wire106[(1'h0):(1'h0)];
  assign wire134 = $unsigned((({(~^wire42), $unsigned(wire109)} ?
                       wire106 : $unsigned(wire109)) ~^ $unsigned(wire43)));
  assign wire135 = $unsigned($unsigned({$unsigned($signed((8'ha8))),
                       $unsigned((^wire133))}));
  assign wire136 = ({$signed(({wire45, wire134} ?
                               {wire108} : wire131[(1'h1):(1'h1)])),
                           ($signed((wire108 <<< wire42)) ?
                               (|$signed(wire41)) : ($unsigned((8'hbd)) && $unsigned(wire109)))} ?
                       $signed(((^~{(8'ha1)}) ?
                           ((-wire86) ?
                               ((8'hae) <= wire110) : {wire135,
                                   (8'hb8)}) : (wire41[(2'h2):(2'h2)] ?
                               $signed(wire43) : (wire134 ?
                                   wire131 : wire108)))) : (&$signed(((~^(7'h43)) >= wire135[(1'h0):(1'h0)]))));
  assign wire137 = ($signed($signed($signed(wire135[(1'h1):(1'h0)]))) | ({$signed($unsigned(wire136))} ?
                       ({(wire133 ? wire110 : wire134)} != ($unsigned(wire109) ?
                           $signed((8'hbf)) : (8'h9f))) : (($unsigned(wire135) ?
                           {(8'hb4)} : (~&wire42)) ^ ($signed(wire45) + (wire131 | wire111)))));
  always
    @(posedge clk) begin
      reg138 <= wire111[(1'h1):(1'h1)];
      reg139 <= wire131[(2'h2):(1'h1)];
      reg140 <= (-$unsigned((^~$signed((wire133 >>> (8'hbe))))));
      if ($unsigned(wire134[(3'h4):(1'h1)]))
        begin
          reg141 <= $signed($unsigned((~&({(8'h9f)} ^~ $unsigned(wire45)))));
          reg142 <= $unsigned(wire111[(4'ha):(3'h5)]);
          if (wire109[(3'h6):(3'h5)])
            begin
              reg143 <= $signed((reg140 ?
                  reg142[(4'hc):(2'h2)] : (~^(~^$unsigned(wire86)))));
              reg144 <= ($unsigned({$signed(reg142[(4'he):(1'h1)])}) ?
                  (($unsigned({wire86, wire133}) - $signed(wire41)) ?
                      wire43 : (|$signed({wire112}))) : ($signed($signed({wire44,
                      wire111})) && (((wire136 ? wire133 : wire134) ?
                      (reg141 ? wire108 : wire135) : (wire111 ?
                          wire86 : wire43)) != $signed(wire43[(3'h4):(3'h4)]))));
            end
          else
            begin
              reg143 <= $signed(wire136[(3'h4):(1'h1)]);
              reg144 <= reg138;
              reg145 <= (!$unsigned(reg138));
              reg146 <= $unsigned(reg141);
            end
          reg147 <= {$signed($unsigned((~^(|wire131)))),
              {(~^$signed(reg145[(3'h6):(3'h4)])),
                  (((~(8'ha0)) ? {reg142} : {wire137, wire131}) - (wire106 ?
                      wire109 : (wire86 > wire133)))}};
          reg148 <= {$unsigned(((wire131[(3'h4):(2'h2)] || ((8'hbd) >> wire45)) ?
                  $unsigned(wire133[(2'h3):(1'h1)]) : $unsigned($signed(wire41))))};
        end
      else
        begin
          reg141 <= ((-reg140) ?
              wire108 : $signed(((^wire42[(4'hc):(3'h6)]) ?
                  $unsigned((~|reg142)) : (&wire45))));
          reg142 <= reg148[(4'hd):(4'hd)];
          reg143 <= ((($unsigned(((8'ha0) ? reg148 : (8'haf))) ?
                      (+reg145) : wire110[(1'h1):(1'h1)]) ?
                  $unsigned($unsigned(((8'hb0) ?
                      wire135 : wire45))) : wire136[(3'h7):(1'h1)]) ?
              ($signed((+(+wire131))) && $signed((8'hb2))) : wire136);
          reg144 <= $signed(reg147[(3'h7):(2'h3)]);
          reg145 <= (!(~|(reg143 ^ $signed((!(8'hae))))));
        end
    end
  assign wire149 = (^~$signed((^~($unsigned((8'haf)) ^ reg139[(2'h2):(1'h1)]))));
  assign wire150 = (-{(~&reg143[(2'h2):(1'h0)])});
  assign wire151 = (!(~^(reg143 >> wire111[(4'hb):(3'h7)])));
  assign wire152 = (~&((+$unsigned($unsigned(wire44))) ? reg143 : wire135));
  assign wire153 = wire136;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module113
#( parameter param129 = ((7'h44) ? (~&(({(8'hac), (8'h9e)} < ((7'h43) ? (8'hb8) : (8'hb6))) != (((7'h43) <= (8'hb5)) ? ((8'hab) ? (8'ha5) : (8'hbe)) : ((8'hbe) < (8'hb2))))) : ({(((8'ha9) ? (8'hbe) : (8'hb1)) ? {(8'hb9)} : ((7'h40) | (8'ha0)))} || ((((8'hbd) == (7'h41)) <= ((8'ha5) >>> (8'hb8))) && (~&(~|(8'hb8))))))
, parameter param130 = (((param129 * (|(~^(8'ha4)))) ? (^~((param129 ? (8'ha2) : param129) >= param129)) : ((-(param129 < (8'h9c))) >= ((^param129) | (~^(8'hba))))) > (param129 ? (((~param129) ? (param129 - param129) : param129) ? ((param129 ? (8'hb7) : (8'ha2)) > (param129 >>> param129)) : {param129, (8'hac)}) : param129)) )
(y, clk, wire117, wire116, wire115, wire114);
  output wire [(32'h81):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h9):(1'h0)] wire117;
  input wire signed [(4'ha):(1'h0)] wire116;
  input wire signed [(3'h7):(1'h0)] wire115;
  input wire [(5'h13):(1'h0)] wire114;
  wire signed [(2'h2):(1'h0)] wire128;
  wire signed [(3'h7):(1'h0)] wire127;
  wire [(4'hd):(1'h0)] wire126;
  wire signed [(5'h11):(1'h0)] wire125;
  wire [(3'h4):(1'h0)] wire124;
  wire [(5'h13):(1'h0)] wire123;
  wire signed [(4'ha):(1'h0)] wire122;
  wire [(4'hb):(1'h0)] wire121;
  wire signed [(5'h14):(1'h0)] wire120;
  wire [(3'h6):(1'h0)] wire119;
  wire signed [(5'h13):(1'h0)] wire118;
  assign y = {wire128,
                 wire127,
                 wire126,
                 wire125,
                 wire124,
                 wire123,
                 wire122,
                 wire121,
                 wire120,
                 wire119,
                 wire118,
                 (1'h0)};
  assign wire118 = wire116[(2'h2):(1'h1)];
  assign wire119 = wire114;
  assign wire120 = (8'ha7);
  assign wire121 = wire120;
  assign wire122 = $unsigned(wire120[(4'hc):(4'hb)]);
  assign wire123 = wire120;
  assign wire124 = ((8'had) << (^~wire120[(5'h14):(4'he)]));
  assign wire125 = (wire120 ?
                       $signed({(+(&wire116)),
                           wire120[(4'hd):(4'hb)]}) : $unsigned((~|{{wire121,
                               wire119}})));
  assign wire126 = ($signed(wire118) ?
                       wire119[(1'h1):(1'h1)] : {(($unsigned(wire116) ?
                               (wire118 ?
                                   wire124 : wire121) : (wire123 >> wire121)) ^ wire125[(5'h11):(4'hd)])});
  assign wire127 = $unsigned($signed($signed(wire122)));
  assign wire128 = ({(~^(wire125 >= (wire114 ? wire127 : wire122)))} ?
                       wire125[(1'h0):(1'h0)] : $unsigned($signed($unsigned((wire116 ^~ wire117)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module88  (y, clk, wire93, wire92, wire91, wire90, wire89);
  output wire [(32'ha0):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h15):(1'h0)] wire93;
  input wire signed [(4'hf):(1'h0)] wire92;
  input wire signed [(4'hc):(1'h0)] wire91;
  input wire signed [(3'h4):(1'h0)] wire90;
  input wire signed [(4'hc):(1'h0)] wire89;
  wire [(5'h11):(1'h0)] wire105;
  wire signed [(4'hc):(1'h0)] wire104;
  wire [(4'hc):(1'h0)] wire103;
  wire [(4'he):(1'h0)] wire102;
  wire signed [(5'h13):(1'h0)] wire101;
  wire [(4'he):(1'h0)] wire100;
  wire [(4'hc):(1'h0)] wire99;
  wire signed [(5'h14):(1'h0)] wire98;
  wire [(4'h8):(1'h0)] wire97;
  wire [(4'he):(1'h0)] wire96;
  wire signed [(4'hb):(1'h0)] wire95;
  wire [(3'h6):(1'h0)] wire94;
  assign y = {wire105,
                 wire104,
                 wire103,
                 wire102,
                 wire101,
                 wire100,
                 wire99,
                 wire98,
                 wire97,
                 wire96,
                 wire95,
                 wire94,
                 (1'h0)};
  assign wire94 = {((!$signed((~wire90))) ?
                          (!(8'hae)) : (-({wire91} ?
                              (wire92 ?
                                  wire90 : wire92) : ((8'hb8) >>> wire91)))),
                      (^((wire93 ^ (wire91 ? wire90 : wire90)) ?
                          $unsigned((8'hb5)) : (|wire92)))};
  assign wire95 = $unsigned($unsigned((((|wire93) << wire92[(3'h6):(3'h6)]) ?
                      wire89[(3'h7):(1'h1)] : wire90[(2'h2):(1'h1)])));
  assign wire96 = (^~{((~(!wire92)) ?
                          $unsigned(((8'ha1) && wire91)) : wire93)});
  assign wire97 = ($unsigned(wire91) ? $signed(wire90[(2'h3):(1'h0)]) : wire93);
  assign wire98 = (^$unsigned(wire89));
  assign wire99 = $signed($signed(((!((8'haa) ^~ (7'h40))) ?
                      wire98[(5'h14):(5'h14)] : ($signed(wire90) * (wire91 >>> wire91)))));
  assign wire100 = (({({wire92} ? $signed((8'hac)) : wire96[(4'hd):(4'hd)])} ?
                       ((wire93[(4'ha):(4'ha)] ?
                           $signed((8'ha3)) : $signed((7'h40))) - $unsigned(wire94)) : wire93) && wire99);
  assign wire101 = $unsigned((&$unsigned($signed((wire92 ? wire99 : wire99)))));
  assign wire102 = ($unsigned({$signed(wire95[(4'hb):(4'h8)])}) ?
                       (wire89 ?
                           wire92[(4'hf):(1'h0)] : $signed(({wire93} | wire99[(3'h7):(3'h7)]))) : ($unsigned((wire89 >>> (wire94 ~^ wire95))) ?
                           ($signed((wire99 != wire93)) ?
                               ((wire97 ? wire90 : wire100) ?
                                   wire91 : ((8'ha0) ?
                                       wire100 : (8'ha0))) : wire92[(4'hd):(3'h4)]) : (8'hb0)));
  assign wire103 = $unsigned(((^~$signed((^wire98))) > ($unsigned((wire95 != wire100)) + $unsigned((wire98 > wire90)))));
  assign wire104 = wire95;
  assign wire105 = {(($signed((wire91 ? wire98 : wire94)) ?
                           $signed($unsigned(wire91)) : ((wire104 >= wire96) << (wire95 ?
                               wire98 : wire97))) << ($unsigned($unsigned((8'h9d))) ?
                           ($unsigned(wire100) ?
                               $unsigned((7'h40)) : $signed(wire95)) : {$unsigned(wire98),
                               wire96[(3'h7):(3'h4)]})),
                       wire97[(4'h8):(1'h0)]};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module46  (y, clk, wire51, wire50, wire49, wire48, wire47);
  output wire [(32'h19d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h2):(1'h0)] wire51;
  input wire [(3'h7):(1'h0)] wire50;
  input wire [(4'ha):(1'h0)] wire49;
  input wire [(5'h10):(1'h0)] wire48;
  input wire [(4'ha):(1'h0)] wire47;
  wire [(4'h9):(1'h0)] wire85;
  wire signed [(5'h10):(1'h0)] wire84;
  reg [(4'hb):(1'h0)] reg83 = (1'h0);
  reg [(4'hc):(1'h0)] reg82 = (1'h0);
  wire [(4'h9):(1'h0)] wire81;
  wire signed [(5'h13):(1'h0)] wire80;
  wire [(2'h2):(1'h0)] wire79;
  wire [(4'h8):(1'h0)] wire78;
  reg [(4'hb):(1'h0)] reg77 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg76 = (1'h0);
  reg [(4'h9):(1'h0)] reg75 = (1'h0);
  reg [(4'h9):(1'h0)] reg74 = (1'h0);
  reg [(5'h15):(1'h0)] reg73 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg72 = (1'h0);
  reg [(2'h3):(1'h0)] reg71 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg70 = (1'h0);
  reg [(4'hc):(1'h0)] reg69 = (1'h0);
  reg [(5'h10):(1'h0)] reg68 = (1'h0);
  reg [(4'he):(1'h0)] reg67 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg66 = (1'h0);
  wire [(4'hd):(1'h0)] wire65;
  wire signed [(5'h15):(1'h0)] wire64;
  wire signed [(5'h11):(1'h0)] wire63;
  wire [(4'ha):(1'h0)] wire62;
  wire signed [(5'h13):(1'h0)] wire61;
  wire signed [(4'h8):(1'h0)] wire60;
  wire signed [(2'h2):(1'h0)] wire59;
  wire [(3'h7):(1'h0)] wire58;
  wire signed [(2'h3):(1'h0)] wire57;
  reg [(5'h12):(1'h0)] reg56 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg55 = (1'h0);
  reg [(4'hf):(1'h0)] reg54 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg53 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire52;
  assign y = {wire85,
                 wire84,
                 reg83,
                 reg82,
                 wire81,
                 wire80,
                 wire79,
                 wire78,
                 reg77,
                 reg76,
                 reg75,
                 reg74,
                 reg73,
                 reg72,
                 reg71,
                 reg70,
                 reg69,
                 reg68,
                 reg67,
                 reg66,
                 wire65,
                 wire64,
                 wire63,
                 wire62,
                 wire61,
                 wire60,
                 wire59,
                 wire58,
                 wire57,
                 reg56,
                 reg55,
                 reg54,
                 reg53,
                 wire52,
                 (1'h0)};
  assign wire52 = ($signed((~^({wire48,
                      wire50} && (wire47 <<< wire50)))) ^ wire50[(2'h2):(2'h2)]);
  always
    @(posedge clk) begin
      reg53 <= (|$signed(wire51));
      reg54 <= wire50;
      reg55 <= reg53[(2'h3):(2'h2)];
      reg56 <= $unsigned((((-(~|wire47)) ?
          wire51[(1'h0):(1'h0)] : (^~reg54)) << (8'hbf)));
    end
  assign wire57 = wire51[(2'h2):(2'h2)];
  assign wire58 = $unsigned((wire51 ?
                      {{$signed(wire52)},
                          ($signed(wire51) ?
                              $unsigned(wire52) : (~wire52))} : (($signed((8'ha1)) ?
                          (!(8'hb9)) : $unsigned(wire51)) <<< wire48[(1'h1):(1'h1)])));
  assign wire59 = $unsigned((~|$signed($signed(wire52))));
  assign wire60 = (!$unsigned($signed((7'h44))));
  assign wire61 = $unsigned({$signed(wire60), (~|wire58)});
  assign wire62 = (wire49[(4'h9):(1'h0)] + wire49[(3'h7):(3'h4)]);
  assign wire63 = $signed(wire49[(3'h4):(1'h0)]);
  assign wire64 = (|($signed($signed((wire51 != (8'ha4)))) ^ (((|wire52) ?
                      wire59 : $unsigned(wire61)) * (+(wire49 ?
                      reg54 : reg56)))));
  assign wire65 = $signed(wire58[(3'h6):(1'h0)]);
  always
    @(posedge clk) begin
      if (wire50[(3'h5):(1'h0)])
        begin
          reg66 <= $unsigned(reg56);
          if ((~&wire52))
            begin
              reg67 <= wire50;
              reg68 <= wire62;
            end
          else
            begin
              reg67 <= wire65[(3'h5):(1'h0)];
              reg68 <= wire61[(3'h4):(2'h2)];
            end
          reg69 <= $signed((($signed((wire61 < wire65)) * $signed((-wire52))) & $signed(wire59[(1'h1):(1'h0)])));
          reg70 <= ((~^((^(reg53 ? wire58 : wire61)) ? reg53 : (^(+wire58)))) ?
              $unsigned($signed($unsigned($unsigned(wire51)))) : {wire63[(2'h2):(1'h1)],
                  (((~^wire62) ?
                      (&(8'hb6)) : (~^wire65)) * (|$unsigned((8'hb1))))});
          if ({$unsigned((8'ha1)), $signed((8'ha3))})
            begin
              reg71 <= $unsigned(((!$signed({reg66, wire58})) ?
                  reg54 : $unsigned(reg68)));
              reg72 <= reg66[(4'hb):(1'h1)];
              reg73 <= wire50;
              reg74 <= $unsigned((&reg72));
              reg75 <= reg53[(2'h3):(2'h2)];
            end
          else
            begin
              reg71 <= ($signed(wire62) ?
                  (|(^~$unsigned(wire63))) : $unsigned((^~((wire59 - (8'hb1)) < (wire51 ?
                      wire51 : reg69)))));
              reg72 <= ((~|$unsigned($unsigned((wire57 | (8'ha1))))) >> $unsigned((|((&wire64) < (reg70 + reg66)))));
              reg73 <= $signed((^({$signed(wire63)} <<< reg74[(1'h1):(1'h1)])));
              reg74 <= $signed(wire65[(1'h1):(1'h1)]);
              reg75 <= wire60[(2'h3):(1'h1)];
            end
        end
      else
        begin
          reg66 <= $unsigned((~((8'ha9) ?
              reg66 : ({wire49} ? wire61 : (wire64 ? reg67 : wire51)))));
          reg67 <= (((|(^reg72[(2'h2):(1'h0)])) || $unsigned(wire50[(2'h3):(1'h1)])) ?
              reg54[(4'ha):(4'h9)] : $unsigned(((~|(8'hae)) ?
                  (~|$unsigned(wire64)) : (~(reg69 > (8'ha1))))));
          reg68 <= (((+($signed(wire64) ? wire51[(1'h1):(1'h1)] : (!wire47))) ?
              ((~&(8'hbe)) != $unsigned(wire59)) : $signed(reg55[(4'hd):(2'h2)])) <<< reg75);
          reg69 <= $signed({$signed((8'hbb))});
        end
      reg76 <= wire64;
      reg77 <= reg53;
    end
  assign wire78 = wire49;
  assign wire79 = reg69;
  assign wire80 = (8'ha7);
  assign wire81 = (-(~|reg76));
  always
    @(posedge clk) begin
      reg82 <= {((+(wire51[(2'h2):(2'h2)] ?
                  $signed(wire48) : (reg70 | reg70))) ?
              {$signed((wire58 ? (8'ha4) : reg73)),
                  ({wire78} <= (^wire57))} : {((wire51 < reg66) || (+(8'haa))),
                  $unsigned(reg76[(1'h0):(1'h0)])}),
          (&(~^reg72[(2'h3):(1'h1)]))};
      reg83 <= $unsigned(({$signed(reg53), wire59} ?
          (^{$signed(wire47)}) : $unsigned($unsigned((wire48 >= reg69)))));
    end
  assign wire84 = (reg66 ?
                      ($unsigned(((reg71 ? wire52 : wire52) ?
                          wire62 : {wire62})) > $unsigned({wire59})) : (+wire60[(3'h4):(2'h2)]));
  assign wire85 = (8'haf);
endmodule