(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h27a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire3;
  input wire signed [(5'h14):(1'h0)] wire2;
  input wire [(5'h14):(1'h0)] wire1;
  input wire signed [(5'h15):(1'h0)] wire0;
  wire [(4'hc):(1'h0)] wire322;
  wire [(5'h14):(1'h0)] wire321;
  reg [(2'h3):(1'h0)] reg320 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg319 = (1'h0);
  reg [(3'h6):(1'h0)] reg318 = (1'h0);
  reg [(3'h4):(1'h0)] reg317 = (1'h0);
  reg [(4'he):(1'h0)] reg316 = (1'h0);
  reg [(4'ha):(1'h0)] reg315 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire314;
  reg signed [(4'hd):(1'h0)] reg313 = (1'h0);
  reg [(5'h12):(1'h0)] reg312 = (1'h0);
  reg signed [(4'he):(1'h0)] reg311 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg310 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg309 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg308 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg307 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg306 = (1'h0);
  reg [(4'he):(1'h0)] reg305 = (1'h0);
  reg [(5'h12):(1'h0)] reg304 = (1'h0);
  wire [(4'hd):(1'h0)] wire303;
  wire [(3'h7):(1'h0)] wire302;
  wire [(2'h3):(1'h0)] wire301;
  wire signed [(4'ha):(1'h0)] wire300;
  reg [(3'h7):(1'h0)] reg299 = (1'h0);
  reg [(5'h11):(1'h0)] reg298 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg297 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg296 = (1'h0);
  reg [(3'h6):(1'h0)] reg295 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg294 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg293 = (1'h0);
  reg [(5'h13):(1'h0)] reg292 = (1'h0);
  reg [(3'h6):(1'h0)] reg291 = (1'h0);
  wire [(5'h13):(1'h0)] wire287;
  wire signed [(4'he):(1'h0)] wire286;
  wire [(4'hb):(1'h0)] wire285;
  wire signed [(4'h9):(1'h0)] wire284;
  wire [(4'h8):(1'h0)] wire283;
  reg signed [(5'h12):(1'h0)] reg282 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg281 = (1'h0);
  reg [(3'h4):(1'h0)] reg280 = (1'h0);
  reg [(4'he):(1'h0)] reg279 = (1'h0);
  reg [(5'h15):(1'h0)] reg278 = (1'h0);
  reg [(5'h15):(1'h0)] reg277 = (1'h0);
  reg [(5'h14):(1'h0)] reg276 = (1'h0);
  reg [(4'hf):(1'h0)] reg275 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg274 = (1'h0);
  reg [(3'h5):(1'h0)] reg273 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg272 = (1'h0);
  wire [(5'h14):(1'h0)] wire271;
  wire signed [(4'he):(1'h0)] wire270;
  wire [(5'h12):(1'h0)] wire269;
  wire signed [(5'h10):(1'h0)] wire268;
  wire [(5'h15):(1'h0)] wire266;
  wire [(2'h3):(1'h0)] wire289;
  assign y = {wire322,
                 wire321,
                 reg320,
                 reg319,
                 reg318,
                 reg317,
                 reg316,
                 reg315,
                 wire314,
                 reg313,
                 reg312,
                 reg311,
                 reg310,
                 reg309,
                 reg308,
                 reg307,
                 reg306,
                 reg305,
                 reg304,
                 wire303,
                 wire302,
                 wire301,
                 wire300,
                 reg299,
                 reg298,
                 reg297,
                 reg296,
                 reg295,
                 reg294,
                 reg293,
                 reg292,
                 reg291,
                 wire287,
                 wire286,
                 wire285,
                 wire284,
                 wire283,
                 reg282,
                 reg281,
                 reg280,
                 reg279,
                 reg278,
                 reg277,
                 reg276,
                 reg275,
                 reg274,
                 reg273,
                 reg272,
                 wire271,
                 wire270,
                 wire269,
                 wire268,
                 wire266,
                 wire289,
                 (1'h0)};
  module4 modinst267 (wire266, clk, wire3, wire1, wire2, wire0, (8'hb0));
  assign wire268 = (($unsigned((wire266[(3'h6):(3'h6)] & $unsigned(wire0))) >>> ((wire1[(4'h8):(3'h5)] ^~ (~(7'h44))) ?
                           ($unsigned(wire0) ^~ $signed(wire1)) : wire266[(3'h4):(1'h1)])) ?
                       {$signed(((wire266 >>> (8'hb5)) <<< {(8'ha2)})),
                           (~^$signed((8'ha7)))} : $signed(((wire266 ?
                           (|wire0) : $signed(wire0)) ^~ {$unsigned(wire266)})));
  assign wire269 = wire0;
  assign wire270 = wire3;
  assign wire271 = ({wire2[(4'hb):(3'h6)],
                           $unsigned((wire269[(3'h4):(2'h3)] + (|wire269)))} ?
                       ((~|$signed($unsigned(wire0))) ?
                           $signed((~(wire1 ?
                               wire3 : (8'hbf)))) : wire270[(2'h3):(1'h1)]) : $unsigned((&{(~wire266),
                           $unsigned((8'ha2))})));
  always
    @(posedge clk) begin
      reg272 <= $signed(($unsigned($unsigned({wire266, wire2})) ?
          (~^$signed(wire1[(4'h9):(1'h0)])) : {{(wire3 > wire271)}}));
      reg273 <= (!{(-{{wire2, wire269}}),
          $unsigned({(~(8'hb4)), (reg272 ? reg272 : wire268)})});
      if ($signed(({wire271[(4'hb):(3'h4)]} ?
          (&wire0[(3'h5):(2'h2)]) : (^~(8'hb0)))))
        begin
          reg274 <= ((!(&($signed(wire269) * (~wire270)))) ?
              $unsigned($unsigned({reg272[(4'h8):(3'h7)]})) : $signed(($signed((&(8'ha8))) || $signed($signed((8'hbb))))));
        end
      else
        begin
          reg274 <= ({(~&($signed((8'hb1)) != wire2[(1'h0):(1'h0)])),
              wire266} * (&(8'h9e)));
          if (reg274[(1'h1):(1'h1)])
            begin
              reg275 <= wire271;
            end
          else
            begin
              reg275 <= {{reg272, (^$unsigned(wire269))}};
              reg276 <= wire1;
              reg277 <= (($signed((wire2[(3'h6):(2'h3)] ^~ $unsigned(wire1))) ?
                  wire2[(4'ha):(4'h8)] : reg274) != $signed(reg276[(2'h3):(2'h2)]));
              reg278 <= (reg274[(2'h2):(1'h1)] ?
                  ($signed(wire3[(3'h6):(2'h3)]) ?
                      ({wire3,
                          $unsigned(reg277)} | $signed(wire2[(4'hb):(4'ha)])) : (~|({reg276} ?
                          reg273[(2'h3):(1'h0)] : $unsigned(wire1)))) : {$signed($signed(wire270))});
            end
          if (wire270[(2'h3):(2'h2)])
            begin
              reg279 <= {(^$unsigned(wire270[(2'h2):(2'h2)]))};
              reg280 <= (((^((reg276 ?
                          (8'h9d) : (8'hb2)) >= reg277[(4'ha):(1'h1)])) ?
                      $signed({reg274[(1'h1):(1'h0)]}) : reg273) ?
                  ($unsigned(((|(8'ha6)) > reg273[(2'h2):(2'h2)])) | wire0) : (-((+((8'hba) ?
                          wire0 : reg273)) ?
                      $unsigned($signed((7'h42))) : ($unsigned(reg276) <= $unsigned((8'hae))))));
              reg281 <= wire2;
            end
          else
            begin
              reg279 <= ($unsigned($unsigned((~$unsigned(wire270)))) ?
                  ($unsigned((&(wire3 || reg275))) ?
                      (^reg276) : ($signed((wire3 ? reg277 : reg278)) ?
                          (+$signed(reg276)) : reg280)) : (reg277[(5'h13):(4'hb)] ?
                      (^(&$signed(reg275))) : ((((8'hb1) ? wire271 : reg279) ?
                              (~^reg280) : (&wire271)) ?
                          reg274 : wire2[(3'h6):(1'h1)])));
              reg280 <= {{$signed($unsigned((reg280 ? (8'ha4) : (8'hbf)))),
                      {$unsigned(wire270)}}};
              reg281 <= wire3[(4'h8):(1'h1)];
              reg282 <= $signed($signed(reg279[(3'h4):(1'h0)]));
            end
        end
    end
  assign wire283 = reg273[(3'h4):(1'h0)];
  assign wire284 = $unsigned(wire0[(1'h0):(1'h0)]);
  assign wire285 = (8'ha7);
  assign wire286 = (wire2 == (wire3 ?
                       (~^$signed(wire1)) : (+(~&$signed(reg276)))));
  module4 modinst288 (.clk(clk), .y(wire287), .wire5(wire0), .wire8(reg276), .wire6(wire266), .wire9(wire268), .wire7(wire284));
  module4 modinst290 (wire289, clk, wire268, wire2, wire1, reg278, reg282);
  always
    @(posedge clk) begin
      if ((wire271[(5'h11):(4'ha)] ?
          $unsigned($unsigned((wire269[(4'hb):(4'ha)] ?
              (reg273 ? (8'hb1) : reg278) : (reg275 ?
                  wire269 : wire1)))) : (($unsigned((reg273 ^ wire283)) ?
                  ($signed((8'ha5)) ?
                      (wire283 | reg282) : wire283[(2'h2):(1'h1)]) : $unsigned($unsigned(reg274))) ?
              $unsigned($signed(wire286[(3'h6):(3'h5)])) : ($unsigned((reg278 ?
                      reg279 : reg276)) ?
                  $unsigned((wire287 ?
                      wire283 : wire0)) : $unsigned((~|wire1))))))
        begin
          reg291 <= (!$signed($signed(wire283[(1'h0):(1'h0)])));
          reg292 <= $signed($unsigned($unsigned($signed(wire289))));
        end
      else
        begin
          reg291 <= reg281;
          reg292 <= {reg272[(2'h2):(1'h0)]};
          reg293 <= (~^((8'hb2) * wire287));
          if ((-{((|$unsigned(wire287)) <= reg282[(4'h8):(2'h2)]),
              {wire3[(4'hc):(1'h0)],
                  {(reg292 ? wire286 : reg273), {wire284, (7'h44)}}}}))
            begin
              reg294 <= wire3;
              reg295 <= (reg291[(1'h0):(1'h0)] <<< (7'h40));
              reg296 <= (~$signed(({$unsigned((8'ha1))} >= (reg273 ?
                  $signed(wire1) : reg282[(1'h0):(1'h0)]))));
            end
          else
            begin
              reg294 <= $unsigned({{(~&$unsigned(reg296)), reg292},
                  (^~wire3[(3'h4):(1'h1)])});
            end
          reg297 <= $signed($signed((+(-((7'h40) ? wire283 : reg294)))));
        end
      reg298 <= {reg276, $signed(reg279[(3'h6):(1'h1)])};
      reg299 <= (+reg272);
    end
  assign wire300 = $signed($signed($signed(reg282)));
  assign wire301 = (!$signed(reg273));
  assign wire302 = (-$unsigned({((wire266 ~^ wire300) >= wire2),
                       (~|$signed(wire266))}));
  assign wire303 = ((|(8'h9d)) ~^ {(((wire1 ? wire283 : reg276) ?
                               (wire283 ? wire285 : wire268) : wire0) ?
                           ($signed(wire284) ~^ (reg297 >= (8'h9f))) : reg272)});
  always
    @(posedge clk) begin
      if (reg275)
        begin
          reg304 <= {wire301, wire303};
          reg305 <= $unsigned(reg272);
          reg306 <= {(^~$unsigned((8'hb5))), wire266};
          if ({(($unsigned((wire289 ? reg304 : reg281)) ?
                      $unsigned((reg304 && wire2)) : reg281[(3'h7):(2'h2)]) ?
                  $signed((^~(^wire284))) : (^((!reg273) ? reg272 : wire285))),
              ($unsigned((~|(wire270 ? reg280 : wire289))) ?
                  reg282 : (reg272[(3'h5):(2'h2)] - (+reg299[(2'h2):(2'h2)])))})
            begin
              reg307 <= $unsigned({reg305});
              reg308 <= $signed($unsigned($unsigned(reg307[(3'h4):(2'h2)])));
              reg309 <= (reg308 ? $signed(wire302) : wire303);
            end
          else
            begin
              reg307 <= ($unsigned(reg293[(3'h4):(1'h0)]) && $signed(wire283[(1'h1):(1'h1)]));
              reg308 <= wire266;
              reg309 <= ($unsigned($unsigned(wire271)) ?
                  ($signed($signed((reg292 < reg304))) - (8'hb6)) : ((8'hb1) + $signed(wire284[(4'h9):(4'h9)])));
            end
          reg310 <= ($unsigned((+((~reg294) ?
              (wire268 - wire285) : (~^reg304)))) + (({wire269,
              {(8'hb7)}} || wire284[(3'h6):(3'h4)]) < wire0[(5'h13):(2'h3)]));
        end
      else
        begin
          reg304 <= ({reg276[(1'h1):(1'h1)]} ?
              (8'ha5) : (reg299[(1'h0):(1'h0)] ?
                  wire283[(3'h7):(1'h1)] : $signed((reg309 ?
                      (wire283 >>> reg276) : (~^wire300)))));
          if ((-{(wire1 ? wire0 : (8'hba))}))
            begin
              reg305 <= {$signed({reg272})};
              reg306 <= (($signed((-wire0)) ?
                      {($signed(wire1) ?
                              (reg293 ?
                                  (8'hb5) : (8'hb7)) : (reg299 >> reg299)),
                          (&(-reg304))} : ((&(reg291 ? reg293 : reg304)) ?
                          reg309 : $signed($unsigned(reg291)))) ?
                  (^~($unsigned((+wire303)) ?
                      wire283[(3'h5):(2'h2)] : reg294)) : {reg306[(2'h2):(2'h2)]});
              reg307 <= $signed($signed((((8'hb9) - wire0) ?
                  wire302[(3'h7):(3'h4)] : wire270[(3'h4):(2'h3)])));
              reg308 <= ((((&wire302) ?
                      reg293 : $signed({reg304})) != (($signed(wire266) << (reg276 <= (8'h9f))) ?
                      wire0 : (~&wire303))) ?
                  (-$unsigned((!(wire3 >> reg304)))) : $unsigned($signed($signed((-reg292)))));
              reg309 <= wire286[(3'h4):(2'h3)];
            end
          else
            begin
              reg305 <= $signed($signed(({$signed(reg297),
                  wire289} != (~&$unsigned(wire3)))));
            end
          reg310 <= wire303;
        end
      reg311 <= $signed(reg274[(5'h10):(4'h8)]);
      reg312 <= reg305;
      reg313 <= reg296;
    end
  assign wire314 = {$unsigned($signed((wire1 ?
                           reg311[(4'ha):(3'h5)] : $unsigned(reg282)))),
                       (-$unsigned(((wire287 >>> reg313) || (&wire287))))};
  always
    @(posedge clk) begin
      if ((~|$signed((^~(|reg282[(1'h1):(1'h1)])))))
        begin
          reg315 <= $unsigned($signed(((&reg312) ?
              $signed((wire270 ?
                  wire268 : wire289)) : (!reg313[(4'hb):(3'h6)]))));
          reg316 <= ($signed((~{(-reg281), reg306})) ?
              reg298 : $signed((wire289 ? (~&reg275) : (|{wire289, (8'hb6)}))));
        end
      else
        begin
          reg315 <= ((({(reg312 || reg278),
                  $signed(wire270)} < $unsigned($signed(wire286))) ?
              $signed($unsigned($unsigned(reg306))) : ((+wire270) ?
                  {$signed(reg278)} : ({reg307} ?
                      reg282[(2'h2):(1'h1)] : reg279[(4'h9):(1'h1)]))) >>> (&$signed($signed($signed(reg315)))));
          if ($signed(((8'ha8) ?
              (($signed(wire284) * $unsigned(wire300)) != (|$signed(reg308))) : {reg279,
                  ($unsigned(reg313) ?
                      $signed(reg305) : (reg279 ? reg281 : (7'h41)))})))
            begin
              reg316 <= wire271;
              reg317 <= ((~wire270) > wire286[(3'h7):(3'h7)]);
            end
          else
            begin
              reg316 <= $signed(reg294[(3'h5):(1'h1)]);
              reg317 <= reg293[(3'h4):(2'h3)];
              reg318 <= ((reg277 ?
                  wire0 : $signed({((8'ha5) & reg281),
                      wire289})) > $signed(reg291));
              reg319 <= (~|$signed($unsigned(reg274)));
            end
        end
      reg320 <= $unsigned(reg293);
    end
  assign wire321 = reg319;
  assign wire322 = reg272;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module4
#( parameter param265 = {((&((&(8'hbe)) - (-(8'h9d)))) ? (^~{((8'haf) < (8'ha9)), ((8'hb8) ? (8'ha4) : (8'hac))}) : (8'ha1)), ((((^(8'ha6)) == ((8'hbb) ? (8'ha6) : (8'ha2))) >>> ({(8'hab), (8'hbf)} >>> (8'h9e))) ? ({((8'h9f) ~^ (7'h42)), ((8'hab) && (8'ha6))} ? (|((8'hbc) ? (8'ha7) : (7'h40))) : ((!(8'ha0)) ? ((8'hbc) ? (8'h9f) : (8'ha1)) : {(8'hba), (8'hbe)})) : ((((8'haa) ? (8'h9f) : (8'hac)) != ((7'h40) < (8'hba))) ? (~^((8'ha1) ^ (8'hb1))) : (^((8'ha7) ^~ (8'hba)))))} )
(y, clk, wire9, wire8, wire7, wire6, wire5);
  output wire [(32'h276):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire9;
  input wire [(5'h14):(1'h0)] wire8;
  input wire signed [(3'h5):(1'h0)] wire7;
  input wire [(5'h15):(1'h0)] wire6;
  input wire [(5'h12):(1'h0)] wire5;
  wire [(4'he):(1'h0)] wire85;
  wire signed [(4'hf):(1'h0)] wire10;
  wire [(2'h2):(1'h0)] wire87;
  wire [(5'h14):(1'h0)] wire88;
  wire [(5'h15):(1'h0)] wire89;
  wire signed [(5'h15):(1'h0)] wire163;
  reg signed [(4'hc):(1'h0)] reg165 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg166 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg167 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg168 = (1'h0);
  reg [(5'h14):(1'h0)] reg169 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg170 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg171 = (1'h0);
  reg [(4'hf):(1'h0)] reg172 = (1'h0);
  reg [(5'h15):(1'h0)] reg173 = (1'h0);
  reg [(5'h10):(1'h0)] reg174 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg175 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg176 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg177 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire178;
  wire [(3'h7):(1'h0)] wire179;
  reg signed [(5'h13):(1'h0)] reg180 = (1'h0);
  reg [(3'h5):(1'h0)] reg181 = (1'h0);
  reg [(4'hf):(1'h0)] reg182 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg183 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg184 = (1'h0);
  reg [(4'he):(1'h0)] reg185 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg186 = (1'h0);
  reg [(4'hc):(1'h0)] reg187 = (1'h0);
  reg [(5'h14):(1'h0)] reg188 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg189 = (1'h0);
  reg [(4'he):(1'h0)] reg190 = (1'h0);
  reg [(5'h14):(1'h0)] reg191 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg192 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg193 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg194 = (1'h0);
  reg [(4'hf):(1'h0)] reg195 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg196 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg197 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire232;
  wire [(4'hd):(1'h0)] wire234;
  reg [(4'h9):(1'h0)] reg235 = (1'h0);
  wire [(5'h11):(1'h0)] wire236;
  wire [(4'h9):(1'h0)] wire237;
  wire [(3'h4):(1'h0)] wire238;
  wire [(5'h13):(1'h0)] wire239;
  wire [(3'h5):(1'h0)] wire240;
  wire [(4'h8):(1'h0)] wire263;
  assign y = {wire85,
                 wire10,
                 wire87,
                 wire88,
                 wire89,
                 wire163,
                 reg165,
                 reg166,
                 reg167,
                 reg168,
                 reg169,
                 reg170,
                 reg171,
                 reg172,
                 reg173,
                 reg174,
                 reg175,
                 reg176,
                 reg177,
                 wire178,
                 wire179,
                 reg180,
                 reg181,
                 reg182,
                 reg183,
                 reg184,
                 reg185,
                 reg186,
                 reg187,
                 reg188,
                 reg189,
                 reg190,
                 reg191,
                 reg192,
                 reg193,
                 reg194,
                 reg195,
                 reg196,
                 reg197,
                 wire232,
                 wire234,
                 reg235,
                 wire236,
                 wire237,
                 wire238,
                 wire239,
                 wire240,
                 wire263,
                 (1'h0)};
  assign wire10 = wire5[(4'he):(4'hd)];
  module11 modinst86 (wire85, clk, wire5, wire7, wire9, wire6, wire10);
  assign wire87 = ($unsigned($unsigned(wire8[(4'h8):(4'h8)])) >> (wire85 ?
                      wire85[(4'hc):(2'h3)] : $unsigned($signed(wire10[(3'h7):(1'h0)]))));
  assign wire88 = (wire9 << $unsigned(wire5[(5'h10):(4'h8)]));
  assign wire89 = $signed(wire9);
  module90 modinst164 (wire163, clk, wire8, wire10, wire89, wire6);
  always
    @(posedge clk) begin
      if ((7'h40))
        begin
          reg165 <= $unsigned($unsigned((^~$signed((wire10 || wire163)))));
          if (wire9[(3'h6):(1'h1)])
            begin
              reg166 <= wire85;
              reg167 <= (($signed(($signed((7'h41)) ?
                      $signed(wire163) : (&wire85))) ?
                  ($unsigned($signed(wire5)) ?
                      wire8[(4'he):(1'h1)] : ($unsigned(wire89) ?
                          (wire85 >= wire163) : (wire87 ?
                              wire89 : wire85))) : (8'hb3)) - $signed((^(~^(~|wire89)))));
            end
          else
            begin
              reg166 <= wire10;
            end
          reg168 <= ((wire89[(5'h10):(4'he)] ?
              (reg165[(1'h1):(1'h0)] ?
                  wire9 : (8'ha2)) : (((~wire9) << $unsigned(wire6)) ^ ((wire6 ?
                      wire89 : (7'h42)) ?
                  reg165 : $signed((8'ha2))))) <<< $unsigned($signed(wire5)));
          reg169 <= $unsigned((((reg168 ? {(8'h9f)} : reg168) > (((8'hbc) ?
                      (8'hae) : wire9) ?
                  $signed(reg168) : $signed((8'hbe)))) ?
              $signed({{wire163}, {wire7}}) : $unsigned($signed((~wire89)))));
          reg170 <= $signed((($signed(wire9[(4'hc):(4'ha)]) ?
              $unsigned((8'ha6)) : wire9[(3'h5):(1'h0)]) < wire87));
        end
      else
        begin
          if (((($unsigned($signed(reg170)) ?
              wire6 : (wire5[(4'hc):(4'h9)] > $unsigned(wire88))) > $signed(wire6[(1'h0):(1'h0)])) != (&$signed($signed($unsigned((8'hbc)))))))
            begin
              reg165 <= ((~|wire8[(4'hb):(3'h5)]) != reg166[(1'h0):(1'h0)]);
              reg166 <= wire163;
              reg167 <= ($signed(wire87) - ($signed(reg165[(4'hc):(4'hc)]) >> ($signed($signed(wire5)) ?
                  wire87[(2'h2):(1'h0)] : $signed({reg170, wire88}))));
              reg168 <= $unsigned(wire9);
            end
          else
            begin
              reg165 <= wire88[(4'h9):(2'h3)];
              reg166 <= (wire89 ?
                  (wire89[(5'h10):(4'hf)] ?
                      (((wire87 + reg165) ?
                          (reg166 ?
                              reg168 : wire9) : ((7'h41) ~^ reg166)) - {wire8,
                          (reg168 <<< wire9)}) : (((wire9 >> wire89) ?
                          $unsigned(reg167) : (~&wire8)) < $unsigned(wire89))) : $signed(((^~(reg170 <<< wire89)) ?
                      $unsigned((wire5 && wire163)) : (~&wire8))));
              reg167 <= ((({(wire85 ? wire9 : reg169)} ?
                      $unsigned($signed(wire9)) : wire87[(1'h1):(1'h1)]) ?
                  wire88[(1'h0):(1'h0)] : $signed(wire89[(3'h6):(2'h3)])) >>> wire163[(5'h15):(5'h11)]);
              reg168 <= wire85;
              reg169 <= $signed($unsigned(($unsigned(wire88[(2'h2):(1'h1)]) ?
                  {(~|wire7)} : {(wire8 ? wire87 : reg167)})));
            end
          reg170 <= (((|($signed(wire7) ?
                  (reg170 ? wire6 : reg168) : $unsigned((8'haa)))) ?
              $signed(wire87) : (~reg169[(5'h11):(4'h9)])) <= wire5);
          if ($signed(($unsigned($signed($unsigned(wire10))) & $signed($signed({reg168,
              wire89})))))
            begin
              reg171 <= reg168;
            end
          else
            begin
              reg171 <= {wire8, (^reg166[(1'h0):(1'h0)])};
              reg172 <= (reg171 ?
                  (wire6 << ($unsigned((~|wire9)) >= wire6[(4'he):(4'hc)])) : reg168[(4'hb):(4'h8)]);
              reg173 <= (-((((reg165 ~^ wire8) & wire89) >= wire9) - $signed($unsigned($signed(reg171)))));
              reg174 <= reg169;
              reg175 <= reg167[(2'h2):(1'h0)];
            end
          reg176 <= $unsigned($signed((+$unsigned((wire8 ? reg166 : wire88)))));
        end
      reg177 <= $signed(reg175);
    end
  assign wire178 = $unsigned(reg172[(2'h3):(1'h1)]);
  assign wire179 = (($signed(wire9) >>> {((wire178 ? reg168 : (8'ha6)) ?
                           (~wire85) : (wire163 <<< reg170))}) == $signed((-((~^(7'h44)) - reg166))));
  always
    @(posedge clk) begin
      reg180 <= ((~|$signed($unsigned(wire163))) ?
          {(wire88 ~^ {(+reg171)}), reg172} : reg169);
      if ({$signed((8'hac)), $unsigned(reg175[(3'h7):(2'h2)])})
        begin
          reg181 <= wire163[(4'he):(4'hc)];
        end
      else
        begin
          if ((({reg174} ? (~$unsigned(reg177)) : (~|reg176)) == reg175))
            begin
              reg181 <= $signed(((wire6[(5'h13):(5'h11)] ?
                  reg180[(5'h12):(4'hf)] : reg174[(1'h1):(1'h0)]) < (^$unsigned($unsigned((8'hb5))))));
              reg182 <= reg165[(4'h9):(3'h6)];
              reg183 <= (reg169 ?
                  (wire5 * wire89) : $unsigned(reg172[(3'h4):(2'h3)]));
              reg184 <= $signed((8'h9d));
              reg185 <= reg173;
            end
          else
            begin
              reg181 <= $signed($unsigned((~&((reg184 || reg167) >= $unsigned(reg171)))));
            end
          reg186 <= reg169;
          reg187 <= {{(wire88[(3'h5):(1'h0)] ? wire87 : (~|(^~reg175)))}};
          if ((+reg185))
            begin
              reg188 <= wire88[(4'hf):(4'ha)];
              reg189 <= reg181;
              reg190 <= wire87[(1'h1):(1'h0)];
              reg191 <= reg172[(4'h9):(1'h1)];
              reg192 <= $unsigned($signed(reg165[(2'h2):(1'h0)]));
            end
          else
            begin
              reg188 <= $signed($signed($unsigned((reg173[(4'hc):(4'hc)] <<< {reg184}))));
              reg189 <= wire178[(4'hb):(3'h6)];
              reg190 <= ($signed($unsigned($unsigned((reg171 << wire7)))) ?
                  ((&($signed(reg188) < reg166)) | {(~$signed(reg188)),
                      wire87}) : ({(reg183 ?
                              $unsigned(reg176) : {(8'haf), reg181})} ?
                      (-wire89) : (~^(~&(wire88 ? wire85 : reg174)))));
              reg191 <= reg180;
            end
        end
      reg193 <= $signed(wire163[(2'h3):(1'h0)]);
      reg194 <= (((7'h43) << (^(8'h9f))) ?
          (8'hb9) : (-$unsigned((reg180 ? $unsigned(reg168) : (&reg170)))));
      reg195 <= $unsigned((wire10 ?
          $unsigned(((^~reg182) * (~wire163))) : (~|(reg190 ?
              $signed(reg168) : $signed((8'h9e))))));
    end
  always
    @(posedge clk) begin
      reg196 <= (reg183[(1'h0):(1'h0)] <<< $signed($unsigned(wire7[(3'h4):(1'h1)])));
      reg197 <= ($unsigned($unsigned(reg188[(5'h11):(5'h10)])) ?
          $unsigned(reg181) : reg177[(3'h6):(2'h3)]);
    end
  module198 modinst233 (.wire199(wire89), .y(wire232), .wire200(reg174), .wire202(reg191), .clk(clk), .wire201(reg193));
  assign wire234 = (reg174 ?
                       (~|reg169) : (wire232[(3'h5):(3'h4)] ?
                           ({(reg185 ? reg188 : wire178),
                               (wire7 ?
                                   reg170 : wire87)} & $unsigned((~&wire89))) : reg194[(2'h2):(2'h2)]));
  always
    @(posedge clk) begin
      reg235 <= (wire9 || (7'h41));
    end
  assign wire236 = (reg192 <= ((wire163 ?
                           reg172[(3'h6):(3'h5)] : reg187[(1'h1):(1'h0)]) ?
                       $unsigned({(reg172 <= wire89), reg171}) : ((~&(8'ha8)) ?
                           ((wire89 ? (8'hba) : wire234) ?
                               (-reg181) : (reg189 ?
                                   reg177 : (8'hba))) : ((wire10 < (8'h9d)) ?
                               (reg183 - reg185) : (reg195 ?
                                   wire7 : wire234)))));
  assign wire237 = ($unsigned($signed($signed($signed(reg176)))) && reg193[(2'h3):(2'h2)]);
  assign wire238 = reg175[(3'h6):(1'h0)];
  assign wire239 = $signed({(reg183 ?
                           (~|reg186) : $signed(reg184[(4'ha):(2'h2)]))});
  assign wire240 = $unsigned((wire89[(5'h14):(5'h14)] ^~ (8'hac)));
  module241 modinst264 (wire263, clk, wire6, wire9, wire8, reg177, reg235);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module241
#( parameter param262 = (&((^~(((8'hb7) ? (8'haa) : (8'hb9)) ? ((8'ha1) <<< (8'ha3)) : {(8'hbc), (8'hbe)})) <= ((~&((8'haa) ? (8'h9c) : (7'h41))) ? (|((8'ha9) ? (7'h43) : (8'h9d))) : (|(^~(8'ha5)))))) )
(y, clk, wire246, wire245, wire244, wire243, wire242);
  output wire [(32'hd1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h2):(1'h0)] wire246;
  input wire signed [(3'h6):(1'h0)] wire245;
  input wire [(3'h4):(1'h0)] wire244;
  input wire [(5'h14):(1'h0)] wire243;
  input wire signed [(3'h6):(1'h0)] wire242;
  reg signed [(5'h13):(1'h0)] reg261 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg260 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg259 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg258 = (1'h0);
  reg [(5'h15):(1'h0)] reg257 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg256 = (1'h0);
  reg [(3'h7):(1'h0)] reg255 = (1'h0);
  reg [(5'h11):(1'h0)] reg254 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg253 = (1'h0);
  reg [(4'hd):(1'h0)] reg252 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire251;
  wire [(3'h4):(1'h0)] wire250;
  wire signed [(5'h15):(1'h0)] wire249;
  wire signed [(4'he):(1'h0)] wire248;
  wire signed [(3'h7):(1'h0)] wire247;
  assign y = {reg261,
                 reg260,
                 reg259,
                 reg258,
                 reg257,
                 reg256,
                 reg255,
                 reg254,
                 reg253,
                 reg252,
                 wire251,
                 wire250,
                 wire249,
                 wire248,
                 wire247,
                 (1'h0)};
  assign wire247 = (-wire244[(2'h3):(1'h0)]);
  assign wire248 = $signed(wire245[(1'h0):(1'h0)]);
  assign wire249 = ($unsigned($signed($signed($unsigned(wire243)))) >>> wire247[(3'h4):(2'h2)]);
  assign wire250 = wire249[(3'h5):(2'h3)];
  assign wire251 = (^~wire246[(1'h0):(1'h0)]);
  always
    @(posedge clk) begin
      if ({$unsigned($unsigned((^wire249[(3'h5):(3'h4)])))})
        begin
          reg252 <= $unsigned(wire242[(1'h1):(1'h1)]);
          reg253 <= (wire247[(1'h1):(1'h1)] ?
              $unsigned($unsigned($signed(wire242))) : ((wire245 ?
                  wire246[(2'h2):(1'h1)] : ((wire249 > wire249) ^~ $signed(wire246))) >> (8'hb9)));
          reg254 <= wire250[(2'h2):(2'h2)];
        end
      else
        begin
          reg252 <= wire245;
          reg253 <= wire250[(3'h4):(3'h4)];
        end
      if (reg253)
        begin
          reg255 <= ({($signed(wire250) ?
                      (8'ha3) : (((8'h9c) ? wire242 : reg253) ?
                          (reg254 ^~ reg253) : (&wire242))),
                  (wire242 ? $unsigned((8'hb4)) : reg253)} ?
              wire246[(1'h1):(1'h1)] : ($unsigned(wire248[(2'h2):(1'h0)]) ?
                  $signed($signed(wire244)) : (reg253 ?
                      (^~(~wire246)) : $unsigned($unsigned(wire249)))));
        end
      else
        begin
          reg255 <= $unsigned(reg255);
          reg256 <= wire250[(1'h0):(1'h0)];
          if ($signed($signed(($unsigned(wire250) ?
              wire250[(2'h3):(1'h0)] : wire243))))
            begin
              reg257 <= ($signed(wire251) <<< reg254[(5'h11):(2'h2)]);
              reg258 <= (wire250[(3'h4):(2'h2)] ?
                  reg252[(3'h6):(3'h4)] : wire245);
              reg259 <= (8'ha5);
              reg260 <= {$signed($unsigned($signed((8'ha7))))};
            end
          else
            begin
              reg257 <= $unsigned(reg256);
              reg258 <= (^~$unsigned(($signed((reg260 >>> reg253)) && $signed({(8'had),
                  wire247}))));
              reg259 <= (!((&$unsigned($unsigned(wire242))) << (($unsigned(wire251) + (reg259 - (8'ha2))) == $signed($signed((8'hb9))))));
            end
          reg261 <= ($signed((reg252 ?
              $unsigned($unsigned(reg259)) : reg256[(4'he):(1'h0)])) <= reg258);
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module198  (y, clk, wire202, wire201, wire200, wire199);
  output wire [(32'h13f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire202;
  input wire signed [(2'h2):(1'h0)] wire201;
  input wire signed [(5'h10):(1'h0)] wire200;
  input wire [(5'h13):(1'h0)] wire199;
  wire [(4'hc):(1'h0)] wire231;
  wire signed [(5'h10):(1'h0)] wire230;
  wire signed [(3'h7):(1'h0)] wire229;
  reg [(4'ha):(1'h0)] reg228 = (1'h0);
  reg [(2'h2):(1'h0)] reg227 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire226;
  reg [(4'hd):(1'h0)] reg225 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg224 = (1'h0);
  reg [(3'h7):(1'h0)] reg223 = (1'h0);
  reg [(5'h13):(1'h0)] reg222 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg221 = (1'h0);
  reg [(2'h2):(1'h0)] reg220 = (1'h0);
  reg [(4'h9):(1'h0)] reg219 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg218 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg217 = (1'h0);
  reg [(2'h3):(1'h0)] reg216 = (1'h0);
  reg [(2'h3):(1'h0)] reg215 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg214 = (1'h0);
  reg [(2'h3):(1'h0)] reg213 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg212 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg211 = (1'h0);
  wire [(4'hf):(1'h0)] wire210;
  wire signed [(4'ha):(1'h0)] wire209;
  reg signed [(5'h12):(1'h0)] reg208 = (1'h0);
  wire [(2'h3):(1'h0)] wire207;
  wire signed [(4'hf):(1'h0)] wire206;
  wire [(4'h8):(1'h0)] wire205;
  reg signed [(5'h10):(1'h0)] reg204 = (1'h0);
  wire [(5'h15):(1'h0)] wire203;
  assign y = {wire231,
                 wire230,
                 wire229,
                 reg228,
                 reg227,
                 wire226,
                 reg225,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 reg219,
                 reg218,
                 reg217,
                 reg216,
                 reg215,
                 reg214,
                 reg213,
                 reg212,
                 reg211,
                 wire210,
                 wire209,
                 reg208,
                 wire207,
                 wire206,
                 wire205,
                 reg204,
                 wire203,
                 (1'h0)};
  assign wire203 = wire199[(2'h2):(1'h0)];
  always
    @(posedge clk) begin
      reg204 <= wire202[(3'h6):(2'h2)];
    end
  assign wire205 = {reg204};
  assign wire206 = wire202;
  assign wire207 = (+{((~&{wire203, wire201}) & wire205), wire205});
  always
    @(posedge clk) begin
      reg208 <= $signed($signed(wire203[(4'hb):(3'h7)]));
    end
  assign wire209 = ({(reg204[(4'h9):(4'h9)] - (wire202 ?
                               $signed((8'hab)) : (&wire201)))} ?
                       (^~$unsigned(wire200)) : reg204);
  assign wire210 = wire199[(5'h12):(2'h2)];
  always
    @(posedge clk) begin
      reg211 <= (((8'haf) ?
          (|((reg208 ? wire203 : wire201) ?
              $unsigned(wire205) : (reg204 ?
                  wire206 : wire209))) : (($signed(wire200) ?
                  wire200[(2'h2):(1'h0)] : $signed(wire199)) ?
              {wire199,
                  $unsigned(wire210)} : wire210[(4'hc):(4'ha)])) && (wire202 << (((|(8'haa)) * {wire206}) ?
          $signed(((8'hb8) ^~ wire201)) : {((8'hbd) ? wire203 : wire201),
              wire205})));
      reg212 <= (8'h9d);
      reg213 <= (~&($unsigned($unsigned((reg204 ?
          wire201 : wire205))) ^~ wire209));
      if (wire205)
        begin
          reg214 <= $unsigned($unsigned($unsigned((~^(|wire209)))));
          if ($unsigned(reg204[(3'h5):(2'h2)]))
            begin
              reg215 <= (^~(-$signed(wire201[(2'h2):(1'h0)])));
              reg216 <= $unsigned($signed(reg212[(1'h0):(1'h0)]));
              reg217 <= reg208[(4'hd):(3'h6)];
              reg218 <= $unsigned($unsigned(reg214[(3'h4):(2'h3)]));
            end
          else
            begin
              reg215 <= $signed(wire201[(1'h1):(1'h1)]);
              reg216 <= (8'ha5);
            end
          reg219 <= ((|$signed(reg204[(3'h7):(3'h6)])) ?
              $signed(wire207) : (($unsigned({reg208, wire205}) ?
                      $signed($unsigned(wire203)) : reg204[(4'hf):(3'h6)]) ?
                  $unsigned(reg213[(1'h0):(1'h0)]) : (~$unsigned((reg211 ?
                      wire210 : (8'ha9))))));
          if ((|$unsigned((^~$unsigned((!wire202))))))
            begin
              reg220 <= {((+$signed(reg212)) > (7'h41))};
              reg221 <= wire199[(4'h9):(2'h3)];
              reg222 <= ((-{(wire207[(2'h2):(1'h0)] ?
                          wire203 : reg204[(4'he):(2'h2)]),
                      (^~$signed((8'ha2)))}) ?
                  $unsigned($signed($signed($signed(wire202)))) : (((^~$unsigned(reg213)) <= $unsigned((8'ha7))) == (^~($signed((8'hb7)) >> $unsigned(wire201)))));
              reg223 <= (reg217[(4'ha):(3'h6)] ?
                  reg219[(2'h3):(1'h0)] : wire201);
            end
          else
            begin
              reg220 <= ($signed((((reg222 ? wire202 : reg223) ?
                      (!reg221) : (reg213 ? reg219 : reg215)) ?
                  $signed((~&wire199)) : ((^reg223) ?
                      (reg216 ^ reg213) : (wire210 ?
                          wire199 : reg216)))) < wire205);
              reg221 <= ({$signed((^(&reg212)))} >>> (8'ha4));
              reg222 <= $signed(wire207);
              reg223 <= (wire209 ?
                  wire201[(1'h0):(1'h0)] : (~&(&$unsigned((reg220 >>> wire205)))));
            end
        end
      else
        begin
          reg214 <= wire200;
          if (wire207)
            begin
              reg215 <= (8'hbf);
              reg216 <= $signed(reg212);
              reg217 <= (({reg217[(4'hc):(4'h8)]} >> (((wire203 <= wire209) ?
                      reg216 : (~|wire203)) ?
                  $unsigned(reg204[(4'h9):(4'h8)]) : (^~$unsigned(reg218)))) < $signed(reg221));
              reg218 <= $signed(reg220);
              reg219 <= (wire203[(5'h15):(4'hc)] << reg223[(1'h1):(1'h1)]);
            end
          else
            begin
              reg215 <= (((8'ha2) ?
                      reg222 : (wire210[(3'h5):(3'h5)] ?
                          (reg223[(3'h4):(2'h2)] && $unsigned(reg220)) : reg204[(1'h0):(1'h0)])) ?
                  reg211 : reg220);
              reg216 <= reg217;
              reg217 <= $unsigned($unsigned(reg215[(1'h0):(1'h0)]));
              reg218 <= wire207[(2'h3):(2'h2)];
            end
          reg220 <= $signed((reg217 ?
              (^wire206[(4'he):(4'h8)]) : reg219[(4'h9):(4'h8)]));
          if ($signed({$signed({$signed(reg223), $signed(reg215)})}))
            begin
              reg221 <= (~^reg213);
            end
          else
            begin
              reg221 <= wire200;
              reg222 <= reg223;
              reg223 <= ($signed(reg211) ?
                  $signed(reg208[(5'h11):(3'h7)]) : $unsigned(wire209));
              reg224 <= (wire202 ?
                  {$signed(((|wire210) ?
                          (wire209 && reg213) : ((8'ha6) ?
                              reg212 : reg212)))} : $unsigned($signed({(wire199 ?
                          wire203 : wire209)})));
            end
          if (reg220)
            begin
              reg225 <= $signed(wire200);
            end
          else
            begin
              reg225 <= (({reg218[(3'h6):(1'h0)]} * $signed(wire209[(1'h1):(1'h1)])) > $signed($signed(reg220[(2'h2):(2'h2)])));
            end
        end
    end
  assign wire226 = reg224;
  always
    @(posedge clk) begin
      reg227 <= ({reg224[(4'hd):(1'h1)]} ?
          $unsigned((^~reg214[(3'h6):(1'h0)])) : {reg213,
              reg218[(3'h7):(1'h1)]});
      reg228 <= (+(~^(~^$unsigned(((8'hb7) ? wire199 : reg222)))));
    end
  assign wire229 = reg212[(2'h2):(2'h2)];
  assign wire230 = (!reg213);
  assign wire231 = ({$signed($signed((wire201 ? wire229 : reg211)))} ~^ reg223);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module90
#( parameter param162 = (&(-({((8'ha0) < (8'hb1))} ? (((8'ha0) ~^ (8'hb8)) ? ((8'hb8) ~^ (8'hab)) : ((8'haf) ^ (8'hb5))) : (((8'ha5) == (8'had)) >> {(8'hbb), (8'hba)})))) )
(y, clk, wire94, wire93, wire92, wire91);
  output wire [(32'h2db):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire94;
  input wire signed [(4'hf):(1'h0)] wire93;
  input wire [(5'h15):(1'h0)] wire92;
  input wire signed [(5'h13):(1'h0)] wire91;
  wire signed [(5'h10):(1'h0)] wire161;
  wire signed [(3'h6):(1'h0)] wire160;
  wire signed [(5'h11):(1'h0)] wire159;
  wire signed [(4'hf):(1'h0)] wire158;
  reg [(5'h15):(1'h0)] reg157 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg156 = (1'h0);
  reg [(5'h13):(1'h0)] reg155 = (1'h0);
  reg signed [(4'he):(1'h0)] reg154 = (1'h0);
  reg signed [(4'he):(1'h0)] reg153 = (1'h0);
  reg [(4'h8):(1'h0)] reg152 = (1'h0);
  reg [(4'hf):(1'h0)] reg151 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg150 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg149 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg148 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg147 = (1'h0);
  reg [(5'h14):(1'h0)] reg146 = (1'h0);
  reg [(3'h7):(1'h0)] reg145 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg144 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg143 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg142 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg141 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg140 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg139 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg138 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg137 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg136 = (1'h0);
  reg [(4'h9):(1'h0)] reg135 = (1'h0);
  reg [(4'hd):(1'h0)] reg134 = (1'h0);
  reg [(4'h8):(1'h0)] reg133 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg132 = (1'h0);
  wire [(4'ha):(1'h0)] wire131;
  reg signed [(3'h7):(1'h0)] reg130 = (1'h0);
  reg [(5'h13):(1'h0)] reg129 = (1'h0);
  reg [(3'h5):(1'h0)] reg128 = (1'h0);
  reg [(5'h13):(1'h0)] reg127 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg126 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg125 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg124 = (1'h0);
  reg [(4'hb):(1'h0)] reg123 = (1'h0);
  reg [(2'h2):(1'h0)] reg122 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg121 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg120 = (1'h0);
  reg [(4'hd):(1'h0)] reg119 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg118 = (1'h0);
  reg [(4'he):(1'h0)] reg117 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg116 = (1'h0);
  reg [(5'h14):(1'h0)] reg115 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg114 = (1'h0);
  reg [(4'hc):(1'h0)] reg113 = (1'h0);
  reg [(3'h5):(1'h0)] reg112 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg111 = (1'h0);
  reg [(4'hd):(1'h0)] reg110 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg109 = (1'h0);
  wire [(3'h5):(1'h0)] wire108;
  wire signed [(4'hb):(1'h0)] wire107;
  wire signed [(5'h13):(1'h0)] wire106;
  reg [(4'h8):(1'h0)] reg105 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg104 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg103 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire102;
  wire [(3'h5):(1'h0)] wire101;
  wire signed [(4'he):(1'h0)] wire100;
  wire [(2'h2):(1'h0)] wire99;
  wire [(3'h6):(1'h0)] wire98;
  wire signed [(4'he):(1'h0)] wire97;
  wire [(2'h3):(1'h0)] wire96;
  wire signed [(4'he):(1'h0)] wire95;
  assign y = {wire161,
                 wire160,
                 wire159,
                 wire158,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 reg149,
                 reg148,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 reg143,
                 reg142,
                 reg141,
                 reg140,
                 reg139,
                 reg138,
                 reg137,
                 reg136,
                 reg135,
                 reg134,
                 reg133,
                 reg132,
                 wire131,
                 reg130,
                 reg129,
                 reg128,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 reg117,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 reg112,
                 reg111,
                 reg110,
                 reg109,
                 wire108,
                 wire107,
                 wire106,
                 reg105,
                 reg104,
                 reg103,
                 wire102,
                 wire101,
                 wire100,
                 wire99,
                 wire98,
                 wire97,
                 wire96,
                 wire95,
                 (1'h0)};
  assign wire95 = ($signed((!(((7'h43) ? wire92 : wire93) ?
                      (7'h43) : (wire94 >>> (7'h41))))) ^~ wire91[(5'h11):(4'he)]);
  assign wire96 = (({$unsigned($unsigned((8'hbc)))} ?
                      (8'hb0) : ((wire94 ^ (|wire92)) ?
                          ($unsigned((8'hbe)) << (wire91 - (8'hb2))) : $unsigned((wire94 ?
                              wire94 : wire95)))) <<< (&(-((wire94 || (8'hb1)) > wire93))));
  assign wire97 = (~|wire94[(1'h1):(1'h0)]);
  assign wire98 = $unsigned((wire95 ?
                      (wire96 * ((wire92 << wire94) ^~ wire97)) : $unsigned(($signed(wire94) ?
                          $unsigned((8'hb6)) : (!wire95)))));
  assign wire99 = ($unsigned((!($unsigned((8'hbe)) ?
                      $unsigned(wire97) : wire97))) ~^ wire94[(4'hf):(2'h3)]);
  assign wire100 = (8'h9c);
  assign wire101 = wire97;
  assign wire102 = $signed(wire99[(2'h2):(1'h0)]);
  always
    @(posedge clk) begin
      reg103 <= wire95;
      reg104 <= (wire99 >= ($signed((wire97 < (~&(8'hbc)))) ?
          (~&$signed(wire102[(1'h0):(1'h0)])) : (wire98 & {(reg103 | (8'hb2)),
              wire92})));
      reg105 <= ((|(reg104 <<< (wire102 || (~&(8'hbc))))) + $unsigned(($unsigned($unsigned(wire94)) ?
          $signed((&wire99)) : (8'hb9))));
    end
  assign wire106 = ({wire99[(1'h0):(1'h0)]} ?
                       $unsigned((!{(|(8'h9f)),
                           {wire98, wire102}})) : (wire92[(4'he):(4'hc)] ?
                           ($unsigned((reg104 ^ wire94)) > wire100) : ((8'hb1) ?
                               wire93 : wire95[(1'h1):(1'h1)])));
  assign wire107 = ($signed($unsigned(wire96)) >>> $signed({reg104,
                       ($signed(wire95) ^ reg105[(2'h2):(1'h0)])}));
  assign wire108 = ({wire106} ~^ (((&$unsigned((8'h9f))) <= (~&((7'h44) <<< (8'ha1)))) > (~|((~|wire92) ?
                       wire107[(3'h7):(3'h4)] : (reg103 ? reg104 : wire101)))));
  always
    @(posedge clk) begin
      if ((((~|wire94[(4'hc):(1'h0)]) <= {wire99[(2'h2):(1'h0)]}) ^~ (8'hb3)))
        begin
          reg109 <= {wire97};
          if ((|$signed($unsigned(((wire98 ? (8'h9d) : wire99) ?
              ((8'hb2) << wire97) : ((8'hb7) * wire100))))))
            begin
              reg110 <= $signed(wire100);
              reg111 <= $signed($signed((wire96 ?
                  wire99 : {wire102[(3'h6):(3'h5)], {wire98}})));
              reg112 <= $unsigned($signed($unsigned(wire92)));
              reg113 <= (wire101 ? reg103 : wire93);
              reg114 <= $unsigned((7'h42));
            end
          else
            begin
              reg110 <= (+wire99);
              reg111 <= wire96;
              reg112 <= (^(|(reg104[(3'h6):(3'h6)] ?
                  wire98[(1'h0):(1'h0)] : $unsigned((^wire95)))));
            end
        end
      else
        begin
          reg109 <= $unsigned({(($signed((8'h9e)) ?
                  reg113[(2'h3):(1'h1)] : (reg112 ?
                      reg105 : (8'haf))) << (-(wire98 ? reg109 : wire108)))});
          reg110 <= (+$signed($signed((reg105[(3'h4):(1'h0)] ?
              (reg114 && wire102) : {wire91}))));
          if ((^~((8'h9f) && (~|{$signed(wire107), (~^wire99)}))))
            begin
              reg111 <= (8'hb8);
              reg112 <= wire96[(2'h3):(1'h1)];
              reg113 <= reg112;
              reg114 <= $unsigned($signed((~{reg105})));
              reg115 <= ((^(&{(wire101 ? wire93 : reg110), (8'ha4)})) ?
                  (~^wire106) : $unsigned($unsigned((^~(wire91 ?
                      reg114 : reg109)))));
            end
          else
            begin
              reg111 <= ((wire94 ?
                      {{(wire98 ? reg113 : wire93)},
                          reg113[(1'h0):(1'h0)]} : ((((7'h42) ?
                              wire97 : wire99) ^~ reg105[(2'h3):(2'h2)]) ?
                          reg111[(2'h3):(2'h2)] : {(wire95 ? wire97 : reg104),
                              (8'hbd)})) ?
                  reg104[(3'h5):(3'h4)] : $signed((^~(~(wire91 ?
                      wire108 : reg111)))));
              reg112 <= $signed({(reg103[(2'h3):(2'h2)] <<< ($signed(wire92) ?
                      $signed(wire98) : ((8'ha1) ? wire93 : reg105))),
                  wire108[(1'h0):(1'h0)]});
              reg113 <= ({$unsigned($signed(wire98)),
                  wire98} == ($signed($unsigned((wire101 >= wire107))) ?
                  (wire97 ?
                      $signed(wire92[(2'h2):(1'h1)]) : ($unsigned(wire106) <<< (8'hab))) : {($signed(wire99) ?
                          (reg109 ? (8'had) : wire101) : ((8'haf) ?
                              reg109 : (8'haf))),
                      wire93}));
            end
        end
      reg116 <= $unsigned((|($signed((reg103 >= wire91)) ?
          wire101 : $signed(reg111[(3'h5):(1'h1)]))));
      reg117 <= $signed({(((|reg105) > (!(8'ha2))) ?
              (+$signed(reg103)) : ((-wire108) >> (reg104 < reg116)))});
    end
  always
    @(posedge clk) begin
      if (reg105[(1'h0):(1'h0)])
        begin
          if (wire100)
            begin
              reg118 <= (~^$unsigned(((8'ha3) ?
                  $signed((wire107 ?
                      reg114 : wire102)) : ($signed(wire99) << (|reg105)))));
              reg119 <= $unsigned({({{reg109, reg117}} ?
                      $unsigned($signed(wire95)) : $unsigned({(8'hb5),
                          wire95}))});
              reg120 <= $signed($signed((^$unsigned(((8'hbd) ?
                  wire106 : wire93)))));
              reg121 <= reg120[(1'h1):(1'h0)];
            end
          else
            begin
              reg118 <= $unsigned({$unsigned($signed({reg105, reg113}))});
              reg119 <= (($unsigned(wire97[(3'h5):(2'h2)]) >>> wire99[(2'h2):(2'h2)]) >> (^~wire107));
            end
          if ({$signed(wire107)})
            begin
              reg122 <= wire99[(1'h0):(1'h0)];
              reg123 <= $unsigned(wire107);
              reg124 <= $signed($signed({reg109[(3'h6):(2'h2)], wire108}));
            end
          else
            begin
              reg122 <= reg121;
              reg123 <= (reg117 | $signed($signed((^~reg115[(4'h9):(1'h1)]))));
              reg124 <= (reg119[(3'h6):(3'h5)] ?
                  wire108[(1'h0):(1'h0)] : {({$signed(reg104)} ?
                          reg103 : reg114[(4'hb):(4'hb)]),
                      (~^$unsigned((reg121 ? reg112 : wire102)))});
            end
          reg125 <= reg105;
          if (($signed((-(^~reg119))) ? (~reg112[(2'h3):(1'h1)]) : reg113))
            begin
              reg126 <= $unsigned(reg103);
              reg127 <= {wire97};
              reg128 <= $signed((!((wire107 ?
                  wire101[(2'h2):(2'h2)] : (reg121 ?
                      reg116 : (8'hb3))) * $unsigned(wire101[(2'h2):(1'h0)]))));
              reg129 <= (|wire107);
            end
          else
            begin
              reg126 <= $signed((~^((~(wire99 >> wire97)) >>> reg112[(3'h4):(1'h0)])));
              reg127 <= {reg126};
              reg128 <= (8'hac);
              reg129 <= $signed((reg126[(3'h7):(2'h2)] ?
                  reg109[(4'h8):(1'h1)] : reg109[(2'h3):(2'h3)]));
              reg130 <= {((~&$unsigned($signed(reg129))) > $unsigned((!reg111[(1'h1):(1'h0)]))),
                  (((|wire101[(1'h1):(1'h1)]) ^ (~&(reg104 ^ wire94))) ?
                      $unsigned($signed((wire98 - reg118))) : (!$signed((~^reg127))))};
            end
        end
      else
        begin
          reg118 <= $signed((8'ha2));
        end
    end
  assign wire131 = $signed($signed(({{(8'ha1), reg104},
                       $unsigned(wire101)} == (reg122[(1'h0):(1'h0)] ?
                       reg110[(3'h4):(1'h0)] : $unsigned((8'ha0))))));
  always
    @(posedge clk) begin
      if (reg124[(3'h4):(3'h4)])
        begin
          reg132 <= (((!(wire96[(2'h2):(2'h2)] >>> wire106)) >>> ((~|$signed(reg123)) * ($signed(reg105) - {(8'ha4)}))) ?
              reg123[(3'h7):(1'h0)] : (~&wire101));
        end
      else
        begin
          if ((reg112 ?
              ($signed($unsigned(reg110[(3'h6):(2'h2)])) * reg103[(2'h2):(1'h0)]) : (-{(+(^~reg127))})))
            begin
              reg132 <= wire106;
              reg133 <= $signed($signed(({$signed((8'hb8)),
                  $unsigned(wire91)} && reg116)));
              reg134 <= ((~&reg122[(1'h1):(1'h1)]) != $signed(reg130[(1'h0):(1'h0)]));
              reg135 <= (~{(8'haa),
                  (((reg129 ? reg104 : reg116) >= reg122) ?
                      ((reg119 ? reg129 : (7'h43)) ?
                          (|(7'h40)) : $unsigned(wire97)) : wire95)});
              reg136 <= (reg115 ?
                  $unsigned(($unsigned((reg112 <= reg112)) == {(reg103 == reg125),
                      reg113[(4'ha):(4'h8)]})) : reg121[(1'h1):(1'h1)]);
            end
          else
            begin
              reg132 <= $unsigned({(!{(reg103 < (8'hb0)), $signed(reg134)}),
                  wire91[(4'hd):(4'hd)]});
              reg133 <= reg135[(3'h7):(2'h2)];
              reg134 <= reg122;
              reg135 <= reg104;
              reg136 <= (-$signed((wire94 ?
                  $unsigned(reg104[(1'h0):(1'h0)]) : (!(+(8'hb9))))));
            end
          if (reg126)
            begin
              reg137 <= wire96[(2'h3):(1'h0)];
              reg138 <= (($unsigned(($unsigned((7'h42)) ?
                      reg129 : (reg111 < wire93))) * (~|(~$unsigned(wire91)))) ?
                  reg128[(1'h1):(1'h1)] : (reg115[(3'h4):(1'h1)] ~^ wire100));
            end
          else
            begin
              reg137 <= (wire97 ?
                  (|$signed(wire91)) : (wire108 ?
                      {($signed(reg138) ? $unsigned(reg137) : reg110),
                          reg104[(3'h7):(2'h3)]} : ($signed($unsigned(wire107)) ?
                          ($signed(reg126) ?
                              (wire94 >>> reg118) : (~|reg128)) : {(~&reg112)})));
              reg138 <= reg120[(4'hb):(3'h7)];
              reg139 <= (~(8'ha7));
              reg140 <= ($signed(reg133) ?
                  (~|$signed(reg114[(4'he):(4'hb)])) : $unsigned({wire97[(4'ha):(3'h4)]}));
              reg141 <= reg140;
            end
        end
      reg142 <= $signed((^$signed($signed($unsigned(reg139)))));
      reg143 <= {{((reg137 + ((8'ha9) ? reg104 : reg109)) ?
                  reg116[(5'h11):(3'h7)] : (~$unsigned(reg132)))}};
      reg144 <= (reg117[(1'h0):(1'h0)] ?
          (|$signed(reg134[(3'h4):(3'h4)])) : reg130[(3'h7):(1'h0)]);
    end
  always
    @(posedge clk) begin
      reg145 <= (&reg123[(3'h4):(2'h3)]);
      reg146 <= $unsigned($signed(reg113));
      if ($signed({(reg134 ?
              $unsigned((|reg114)) : $unsigned($unsigned(reg136))),
          $unsigned($signed((wire92 ^ wire95)))}))
        begin
          reg147 <= $signed({reg113});
          reg148 <= ((^~(8'haf)) ? $signed(reg103) : reg128);
          if (($signed($unsigned($signed(wire98[(3'h5):(1'h1)]))) - (($signed((reg135 <<< wire97)) >>> $signed(reg124[(1'h0):(1'h0)])) > $unsigned($unsigned((reg129 ~^ reg123))))))
            begin
              reg149 <= $signed((|$signed(reg142[(3'h6):(3'h5)])));
            end
          else
            begin
              reg149 <= $unsigned($signed($unsigned((wire93[(3'h7):(3'h5)] >>> reg133))));
            end
          reg150 <= (^~((+(8'hbf)) ? wire98 : $signed((|$unsigned((7'h42))))));
          reg151 <= $signed((^~$signed($unsigned(reg136))));
        end
      else
        begin
          reg147 <= ($unsigned((!(~|$signed((8'ha9))))) && $signed({($unsigned((8'hba)) ?
                  (reg115 ? wire101 : (8'hba)) : (wire100 == reg146))}));
          reg148 <= ($unsigned($signed($signed((8'hb1)))) ?
              (~&$signed(({reg127,
                  reg134} << reg126))) : (+$signed(reg126[(2'h3):(2'h2)])));
          reg149 <= ({$unsigned(((reg147 * (8'hbb)) ?
                      (reg134 * (8'hab)) : {wire107, reg148})),
                  reg147[(2'h2):(1'h1)]} ?
              $signed(({$unsigned(reg118)} << (reg135 & reg117[(3'h4):(1'h1)]))) : ((+(8'ha0)) ^~ {($unsigned(reg125) <= (!reg140))}));
          reg150 <= ($signed((($unsigned((8'hb0)) || reg141) ?
                  (^~reg112[(2'h2):(2'h2)]) : reg123)) ?
              (~&reg113) : ($signed($unsigned($unsigned(reg123))) ?
                  $unsigned(((reg103 ?
                      reg117 : reg130) <= $unsigned((7'h43)))) : ((reg128[(2'h2):(2'h2)] ?
                          wire108 : wire108[(3'h4):(3'h4)]) ?
                      $unsigned(wire108) : ($unsigned(reg130) ?
                          reg105 : (reg134 == reg112)))));
        end
      if (reg110)
        begin
          if (((reg118 ?
                  $unsigned((^~(~^reg134))) : $signed(($unsigned(reg145) ?
                      {wire106} : reg129))) ?
              reg147[(3'h6):(3'h4)] : (~(^{reg110[(4'h9):(1'h1)]}))))
            begin
              reg152 <= reg120[(3'h6):(2'h2)];
            end
          else
            begin
              reg152 <= (~&$unsigned(reg149));
              reg153 <= $unsigned(wire96);
              reg154 <= ($signed(($unsigned((wire107 ?
                  wire96 : reg152)) || {reg150,
                  (reg145 * reg147)})) && $signed({(((8'h9d) ?
                      reg127 : reg149) <= reg130),
                  $signed(reg125[(4'ha):(3'h4)])}));
              reg155 <= $signed({$unsigned((&(reg105 ? (8'hb3) : reg150))),
                  $unsigned(((8'h9f) & (!wire96)))});
            end
          reg156 <= reg133;
          reg157 <= ((+(!({reg156} & $signed(reg153)))) ?
              {wire107[(2'h3):(2'h2)],
                  (~&((wire91 ? reg135 : reg120) ?
                      $unsigned(wire92) : {reg142}))} : ($signed(reg152[(4'h8):(3'h6)]) ^~ $unsigned((reg136 + (reg144 && reg103)))));
        end
      else
        begin
          reg152 <= $unsigned(reg151);
          reg153 <= $unsigned(({wire108} ?
              (|(8'ha5)) : (^((reg133 ? reg118 : wire131) ?
                  {reg143} : (reg119 ? reg115 : reg141)))));
          reg154 <= (&(|reg146[(3'h7):(3'h6)]));
        end
    end
  assign wire158 = (($signed((~^(reg141 | reg144))) ?
                           (8'ha1) : reg152[(2'h3):(1'h0)]) ?
                       $signed((reg150[(3'h7):(2'h2)] >>> {$unsigned((8'hb6)),
                           reg157[(4'h9):(2'h2)]})) : reg104[(3'h5):(1'h0)]);
  assign wire159 = reg132;
  assign wire160 = (((~|{$unsigned(reg146)}) ?
                       $unsigned($unsigned(reg154)) : ($signed((reg152 != reg149)) - ((^(7'h43)) >> (reg125 * (8'had))))) + (((|reg115) ~^ $unsigned($signed(wire98))) != reg121[(1'h1):(1'h0)]));
  assign wire161 = (((~(~^reg118[(2'h3):(2'h3)])) >= wire93[(3'h7):(3'h5)]) ?
                       (~(~|(reg103 << reg146))) : (reg123[(2'h3):(1'h0)] ?
                           reg141 : (^~(^(8'hbf)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module11  (y, clk, wire16, wire15, wire14, wire13, wire12);
  output wire [(32'h31e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h8):(1'h0)] wire16;
  input wire signed [(3'h4):(1'h0)] wire15;
  input wire signed [(4'hc):(1'h0)] wire14;
  input wire signed [(4'hf):(1'h0)] wire13;
  input wire signed [(3'h7):(1'h0)] wire12;
  reg signed [(2'h3):(1'h0)] reg84 = (1'h0);
  reg [(4'ha):(1'h0)] reg83 = (1'h0);
  reg [(5'h12):(1'h0)] reg82 = (1'h0);
  reg [(4'he):(1'h0)] reg81 = (1'h0);
  reg [(4'hc):(1'h0)] reg80 = (1'h0);
  reg [(2'h2):(1'h0)] reg79 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg78 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg77 = (1'h0);
  reg [(5'h15):(1'h0)] reg76 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg75 = (1'h0);
  reg [(2'h3):(1'h0)] reg74 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg73 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg72 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg71 = (1'h0);
  reg [(5'h14):(1'h0)] reg70 = (1'h0);
  reg [(3'h6):(1'h0)] reg69 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg68 = (1'h0);
  reg [(4'h8):(1'h0)] reg67 = (1'h0);
  reg [(3'h6):(1'h0)] reg66 = (1'h0);
  reg [(5'h10):(1'h0)] reg65 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg64 = (1'h0);
  reg [(4'he):(1'h0)] reg63 = (1'h0);
  reg [(3'h6):(1'h0)] reg62 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg61 = (1'h0);
  reg [(5'h13):(1'h0)] reg60 = (1'h0);
  reg [(3'h7):(1'h0)] reg59 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg58 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg57 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg56 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg55 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg54 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg53 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg52 = (1'h0);
  reg [(3'h5):(1'h0)] reg51 = (1'h0);
  reg [(3'h6):(1'h0)] reg50 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg49 = (1'h0);
  reg [(3'h5):(1'h0)] reg48 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg47 = (1'h0);
  reg [(5'h11):(1'h0)] reg46 = (1'h0);
  reg signed [(4'he):(1'h0)] reg45 = (1'h0);
  reg signed [(4'he):(1'h0)] reg44 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg43 = (1'h0);
  reg [(4'hc):(1'h0)] reg42 = (1'h0);
  reg [(5'h15):(1'h0)] reg41 = (1'h0);
  reg [(4'h8):(1'h0)] reg40 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg39 = (1'h0);
  wire [(4'he):(1'h0)] wire38;
  wire [(5'h15):(1'h0)] wire37;
  wire [(5'h10):(1'h0)] wire36;
  wire [(3'h7):(1'h0)] wire35;
  wire [(4'hd):(1'h0)] wire34;
  reg [(4'hf):(1'h0)] reg33 = (1'h0);
  wire [(5'h11):(1'h0)] wire32;
  wire signed [(4'hb):(1'h0)] wire31;
  wire signed [(5'h10):(1'h0)] wire30;
  reg [(5'h12):(1'h0)] reg29 = (1'h0);
  reg [(3'h4):(1'h0)] reg28 = (1'h0);
  reg [(4'he):(1'h0)] reg27 = (1'h0);
  reg [(4'hd):(1'h0)] reg26 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg25 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg24 = (1'h0);
  reg [(5'h11):(1'h0)] reg23 = (1'h0);
  reg [(3'h4):(1'h0)] reg22 = (1'h0);
  wire [(2'h3):(1'h0)] wire21;
  wire [(4'hc):(1'h0)] wire20;
  wire [(4'h8):(1'h0)] wire19;
  wire [(5'h15):(1'h0)] wire18;
  wire signed [(3'h6):(1'h0)] wire17;
  assign y = {reg84,
                 reg83,
                 reg82,
                 reg81,
                 reg80,
                 reg79,
                 reg78,
                 reg77,
                 reg76,
                 reg75,
                 reg74,
                 reg73,
                 reg72,
                 reg71,
                 reg70,
                 reg69,
                 reg68,
                 reg67,
                 reg66,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 reg55,
                 reg54,
                 reg53,
                 reg52,
                 reg51,
                 reg50,
                 reg49,
                 reg48,
                 reg47,
                 reg46,
                 reg45,
                 reg44,
                 reg43,
                 reg42,
                 reg41,
                 reg40,
                 reg39,
                 wire38,
                 wire37,
                 wire36,
                 wire35,
                 wire34,
                 reg33,
                 wire32,
                 wire31,
                 wire30,
                 reg29,
                 reg28,
                 reg27,
                 reg26,
                 reg25,
                 reg24,
                 reg23,
                 reg22,
                 wire21,
                 wire20,
                 wire19,
                 wire18,
                 wire17,
                 (1'h0)};
  assign wire17 = (!{wire12, (|(|$unsigned((8'hb6))))});
  assign wire18 = (^~(|$signed((|(wire17 != wire12)))));
  assign wire19 = (~|wire12);
  assign wire20 = ({$unsigned(((8'hba) ?
                          $unsigned(wire15) : wire17[(3'h5):(2'h3)]))} >> (wire17 > (|$signed($signed(wire18)))));
  assign wire21 = ($unsigned($unsigned(((wire14 > wire18) ?
                      $unsigned((7'h44)) : (~&wire18)))) * (wire18[(4'hc):(3'h5)] ?
                      wire15 : wire18));
  always
    @(posedge clk) begin
      reg22 <= ({$unsigned($signed($signed(wire13)))} ^~ $signed($unsigned({(|wire19),
          ((7'h40) << wire21)})));
      reg23 <= (wire17 > {$unsigned((-(wire15 >= wire20))),
          ((^$unsigned(wire18)) ?
              (wire12[(1'h0):(1'h0)] ?
                  (~wire15) : (wire14 == wire13)) : (((8'ha2) ?
                  wire16 : wire14) <<< $signed(wire14)))});
      reg24 <= (&reg23[(4'hd):(4'hc)]);
      if (reg23)
        begin
          reg25 <= $unsigned($signed((8'hac)));
        end
      else
        begin
          if ((wire13[(4'hf):(4'ha)] ^~ $signed($unsigned((~{wire19})))))
            begin
              reg25 <= wire12;
            end
          else
            begin
              reg25 <= (+($signed($signed($signed(wire18))) ?
                  (((wire17 << (8'ha0)) >= $signed(reg22)) >>> {(^~wire12)}) : $unsigned(((reg23 ?
                          reg25 : wire13) ?
                      $unsigned(wire19) : reg22))));
              reg26 <= ($unsigned(($signed({wire20}) ?
                      wire16[(2'h2):(2'h2)] : {$signed((8'ha4))})) ?
                  (-$signed((8'haf))) : ($signed(wire14[(4'h8):(4'h8)]) & wire15));
            end
          reg27 <= {(~|(wire18 ?
                  $unsigned($unsigned(wire17)) : $unsigned((wire16 ?
                      (7'h40) : reg24)))),
              ($signed((+$unsigned(wire13))) ?
                  $unsigned($unsigned((^wire21))) : (~^wire20[(4'h8):(3'h6)]))};
          reg28 <= {wire12};
        end
      reg29 <= (^$unsigned((({wire12, reg22} || reg27) < $unsigned(wire12))));
    end
  assign wire30 = wire12;
  assign wire31 = reg22;
  assign wire32 = $signed(wire16[(3'h5):(2'h2)]);
  always
    @(posedge clk) begin
      reg33 <= (^(~^$unsigned(wire32[(4'h9):(3'h7)])));
    end
  assign wire34 = {(((-(^reg28)) ^~ (+(wire32 ? reg25 : (8'hbc)))) ?
                          (8'hb4) : wire31)};
  assign wire35 = (reg22[(1'h1):(1'h0)] ?
                      wire18 : {($signed(wire13[(3'h7):(2'h3)]) ?
                              (~|$signed(wire18)) : wire13[(1'h0):(1'h0)]),
                          $unsigned(reg22)});
  assign wire36 = wire19;
  assign wire37 = $signed($unsigned((~&wire19[(3'h5):(2'h3)])));
  assign wire38 = reg22[(2'h2):(1'h0)];
  always
    @(posedge clk) begin
      reg39 <= reg28;
      if (reg27[(4'he):(4'he)])
        begin
          reg40 <= ($signed(wire16[(3'h5):(3'h4)]) + {({$unsigned(reg33),
                  reg39[(5'h10):(2'h2)]} < reg22)});
          reg41 <= (^{(~|$unsigned($unsigned(reg39)))});
          reg42 <= wire16[(1'h1):(1'h0)];
          reg43 <= reg29;
          reg44 <= wire34;
        end
      else
        begin
          reg40 <= $signed($unsigned((((wire21 + wire13) ? (!reg43) : wire34) ?
              $signed($signed(reg40)) : ((reg44 < wire31) ?
                  $signed(wire37) : (reg22 <= wire20)))));
          reg41 <= reg43[(4'h8):(4'h8)];
          reg42 <= (^reg41);
          reg43 <= $signed(($unsigned($unsigned((wire21 ?
              wire15 : reg23))) >>> (~|(~^((8'hb1) ^~ wire17)))));
        end
      reg45 <= (wire34[(4'h8):(3'h5)] ?
          $unsigned(wire36[(4'h9):(2'h3)]) : (~(~|($signed(reg33) ?
              (^~(8'hb2)) : $unsigned(wire30)))));
      reg46 <= (+reg33[(4'h9):(2'h2)]);
    end
  always
    @(posedge clk) begin
      reg47 <= (({wire15[(1'h0):(1'h0)], (8'hbe)} ?
          reg26[(3'h5):(2'h2)] : (^(^~wire19))) ^~ ((8'hbd) <<< {wire32[(1'h0):(1'h0)],
          (~|$signed(wire18))}));
      reg48 <= (reg43 + ($signed((reg22 - ((7'h40) > reg46))) != (-({reg41} && (&wire12)))));
      if ($signed((8'hba)))
        begin
          reg49 <= ($signed((reg28 * (-(reg39 ?
              wire16 : wire35)))) >>> (wire32[(4'hb):(3'h5)] + $unsigned(((reg23 | reg41) ?
              reg48 : reg29[(5'h11):(3'h6)]))));
          if ((wire35[(3'h5):(3'h5)] * $unsigned(reg28)))
            begin
              reg50 <= wire36;
              reg51 <= wire32;
              reg52 <= (~&$signed((8'hb2)));
              reg53 <= {(reg27 ? wire34[(1'h1):(1'h1)] : reg40[(3'h6):(1'h1)])};
            end
          else
            begin
              reg50 <= (wire17 << wire15);
              reg51 <= (wire31 ?
                  $unsigned((($unsigned(reg43) ? reg28 : (wire15 ~^ wire17)) ?
                      $signed((^reg22)) : wire30)) : $signed((&$signed((~^(7'h40))))));
            end
          reg54 <= $signed(reg49);
          reg55 <= $unsigned(($unsigned(($signed(wire38) ?
                  $signed(wire37) : ((8'hb6) >>> wire32))) ?
              reg50 : $signed(((&wire35) ?
                  wire35[(3'h5):(1'h1)] : (wire14 || wire32)))));
        end
      else
        begin
          reg49 <= (!($unsigned(reg23[(3'h7):(1'h1)]) ?
              $signed((reg55 ?
                  $signed(reg42) : wire20)) : ($signed($unsigned(reg27)) ?
                  wire12 : (((7'h40) ? reg44 : wire20) && $unsigned(wire12)))));
          if (reg40)
            begin
              reg50 <= $signed(reg22);
              reg51 <= {wire34,
                  $signed(($unsigned($signed(wire21)) ?
                      (8'h9d) : $unsigned((reg23 ? reg52 : wire15))))};
              reg52 <= ($signed(((reg48 ?
                      (wire32 && wire34) : $signed(wire32)) >= reg45[(1'h1):(1'h1)])) ?
                  wire12[(3'h4):(3'h4)] : (~reg40));
              reg53 <= (!reg43);
            end
          else
            begin
              reg50 <= {reg52, reg48[(2'h3):(2'h2)]};
            end
          reg54 <= (|(|(^~(~^wire34))));
        end
    end
  always
    @(posedge clk) begin
      reg56 <= (wire32 ? reg33[(2'h3):(2'h3)] : wire31[(1'h1):(1'h1)]);
      if (reg48)
        begin
          reg57 <= (-reg51[(3'h4):(1'h0)]);
          reg58 <= (8'hb1);
          reg59 <= ((&reg29[(4'h8):(2'h3)]) | {($signed({(8'hb4)}) ?
                  reg41[(5'h11):(5'h10)] : $signed(reg45))});
          reg60 <= ($unsigned($unsigned((^~(!wire20)))) ?
              $unsigned($unsigned((+$signed(reg52)))) : reg39);
        end
      else
        begin
          reg57 <= (((reg51[(1'h1):(1'h1)] ?
                      (~&((8'hbc) ?
                          reg50 : reg54)) : $unsigned(reg55[(4'h9):(4'h8)])) ?
                  reg44[(1'h1):(1'h0)] : {reg59, (|reg26)}) ?
              reg29[(3'h5):(3'h5)] : $signed(((!$signed((8'h9e))) ~^ reg54[(3'h7):(2'h3)])));
          reg58 <= ((8'hb2) >= reg50[(2'h2):(1'h0)]);
          reg59 <= reg23;
          reg60 <= $unsigned((|(8'h9e)));
        end
      if ($unsigned($unsigned(wire20[(1'h1):(1'h0)])))
        begin
          if (wire35[(2'h2):(1'h0)])
            begin
              reg61 <= reg44[(1'h0):(1'h0)];
              reg62 <= ((reg22 ?
                  reg57[(1'h0):(1'h0)] : reg24) == $signed(({$signed(reg22),
                  (wire30 ? reg39 : reg48)} != $signed(((7'h42) | wire12)))));
              reg63 <= reg44;
              reg64 <= $signed({$unsigned(reg53[(4'h9):(3'h6)])});
              reg65 <= (~|$unsigned(((reg47 ?
                  $unsigned(reg55) : (~reg51)) ~^ $signed(reg51[(2'h3):(2'h3)]))));
            end
          else
            begin
              reg61 <= reg58;
              reg62 <= (-reg26);
            end
          reg66 <= (reg50[(2'h3):(1'h1)] <= ({(^$unsigned((8'hb3)))} <= reg22[(1'h1):(1'h0)]));
          if ({$unsigned(reg41)})
            begin
              reg67 <= ((((~&reg52) ?
                      ((^reg66) >> $unsigned(wire32)) : {$signed(reg28),
                          $unsigned(reg39)}) ?
                  $signed((~^{reg47,
                      (7'h42)})) : $unsigned(({wire12} << $signed(reg43)))) ^~ (((|(reg60 - reg50)) ?
                  reg39[(4'hb):(4'h9)] : reg45) * ({(wire15 ^ reg51),
                  $unsigned(reg27)} - $unsigned(wire32))));
              reg68 <= (~((($signed(reg53) * (8'ha7)) ^ {reg49[(2'h3):(2'h2)]}) >>> reg48));
              reg69 <= $signed(wire31[(3'h5):(3'h4)]);
              reg70 <= ((({(wire15 ? reg47 : reg53)} ?
                          ((8'hb9) ?
                              $unsigned((8'hb7)) : {(7'h43), reg57}) : wire18) ?
                      $unsigned(($unsigned(reg33) <= (reg68 || wire31))) : $unsigned($unsigned({reg52}))) ?
                  reg61 : reg54[(3'h4):(3'h4)]);
              reg71 <= reg45[(4'h9):(1'h0)];
            end
          else
            begin
              reg67 <= (({({reg29, reg23} ?
                          $unsigned((8'hb7)) : {(8'ha3), (8'hb8)})} ?
                  $unsigned((wire14 ?
                      wire21 : ((8'hba) ?
                          (8'hbb) : reg39))) : $unsigned($unsigned(reg71))) + ((~|reg57) ?
                  (reg61[(4'hd):(4'h8)] ?
                      $unsigned(((8'hbe) ?
                          reg25 : wire35)) : $signed($signed(wire38))) : ((reg46[(4'he):(3'h7)] ?
                          (reg71 - reg65) : $signed(wire20)) ?
                      {(wire35 ^~ reg47)} : ((~&wire15) ?
                          $signed(reg54) : $unsigned(reg27)))));
              reg68 <= (reg27 <<< $unsigned({(|(reg24 ? wire18 : (8'ha3)))}));
              reg69 <= $signed($unsigned($signed($signed($unsigned(reg40)))));
            end
          if (reg28[(3'h4):(3'h4)])
            begin
              reg72 <= (~^(^(($unsigned(wire38) * wire30[(2'h3):(2'h3)]) ?
                  $unsigned(wire36[(4'hd):(1'h0)]) : ($signed(reg70) << (reg71 & reg59)))));
              reg73 <= wire16;
              reg74 <= (($signed($unsigned((~|reg48))) ?
                      ($unsigned((wire38 ? reg25 : reg46)) ~^ $unsigned((reg45 ?
                          reg23 : reg48))) : wire34) ?
                  reg54 : {wire17[(3'h5):(2'h3)]});
              reg75 <= ($unsigned(reg65) != (reg33[(2'h2):(1'h0)] ?
                  reg66[(1'h0):(1'h0)] : (8'hb7)));
              reg76 <= reg45;
            end
          else
            begin
              reg72 <= $signed(reg39[(4'h8):(2'h2)]);
              reg73 <= $unsigned($unsigned(((~|{(8'ha4)}) <<< {(reg45 ?
                      reg39 : reg76)})));
              reg74 <= reg76;
              reg75 <= reg75;
              reg76 <= (&$signed({(reg28[(3'h4):(2'h3)] ?
                      {wire30} : (^reg48))}));
            end
        end
      else
        begin
          reg61 <= (~|{$unsigned(((7'h42) <= reg25[(1'h0):(1'h0)])),
              reg25[(1'h0):(1'h0)]});
        end
      if (($signed(($signed(reg41) * reg63[(2'h3):(2'h2)])) <= ((reg26 - reg63[(4'hd):(4'h9)]) <<< (reg41 ~^ ({reg50} * ((7'h42) ?
          reg23 : (8'ha5)))))))
        begin
          reg77 <= reg59;
          reg78 <= (wire14[(4'hc):(4'ha)] <= $signed($signed($signed((wire35 == reg52)))));
          reg79 <= {((($signed(reg55) ?
                      (reg76 ?
                          reg68 : wire31) : (reg41 * wire15)) < $unsigned(reg44[(4'h8):(1'h1)])) ?
                  ({reg61, $unsigned(wire15)} ?
                      (!(!reg58)) : $signed(reg48[(2'h3):(2'h2)])) : (!$unsigned($unsigned(wire20))))};
          if (reg69[(3'h4):(1'h0)])
            begin
              reg80 <= (reg44[(3'h6):(1'h0)] ?
                  (wire34 ?
                      reg40 : $signed(reg72[(3'h7):(3'h4)])) : (~&$unsigned($signed((~|reg47)))));
              reg81 <= wire16;
              reg82 <= (~|reg47);
            end
          else
            begin
              reg80 <= reg49[(3'h4):(3'h4)];
              reg81 <= wire31;
            end
        end
      else
        begin
          if ((8'h9f))
            begin
              reg77 <= ($signed(({(~^reg59)} | $signed((reg47 ~^ wire16)))) >> (|(^~reg25)));
              reg78 <= ($unsigned((reg61[(3'h5):(1'h1)] == ($signed(reg28) ?
                  reg67 : ((8'hb2) ?
                      wire30 : wire21)))) <<< (reg67 ^ $signed($unsigned(reg25[(3'h4):(2'h3)]))));
              reg79 <= ($unsigned(reg22) ?
                  $unsigned(reg80) : (~^{wire16[(2'h2):(2'h2)],
                      $unsigned(reg53)}));
            end
          else
            begin
              reg77 <= (reg68 * $unsigned(wire35));
              reg78 <= reg39[(4'h8):(3'h7)];
            end
          if ((~{$signed((7'h44)),
              ({reg82[(4'hd):(4'hb)]} | {$signed(reg80)})}))
            begin
              reg80 <= ($signed((((reg46 ^~ reg80) ~^ reg75) >> wire21)) ~^ $unsigned(((~&$unsigned(wire19)) << $signed($signed((8'hbf))))));
              reg81 <= {{{$signed((|reg79)), $unsigned(reg63)}},
                  $signed(wire37[(3'h5):(1'h1)])};
              reg82 <= (reg71[(2'h2):(1'h0)] ?
                  $signed($unsigned($signed($signed(wire14)))) : reg22[(1'h1):(1'h1)]);
              reg83 <= $unsigned($signed(((^~(+reg46)) ?
                  $unsigned((wire30 ? reg68 : wire34)) : {wire15,
                      reg60[(1'h0):(1'h0)]})));
              reg84 <= ((reg65 <<< (+((+reg70) >>> wire15))) ?
                  $unsigned({reg43[(4'h8):(3'h4)]}) : $unsigned((reg72[(1'h0):(1'h0)] ?
                      $unsigned({wire31, wire17}) : {{reg71, reg50}, reg73})));
            end
          else
            begin
              reg80 <= (($unsigned($unsigned((7'h41))) ?
                  $unsigned($unsigned((~reg40))) : (7'h41)) || (^~(($signed(reg23) ?
                      (8'hbf) : wire37[(4'hc):(4'h8)]) ?
                  wire17[(3'h5):(2'h3)] : (^~((8'ha3) || reg62)))));
              reg81 <= (($signed({(|reg80)}) ?
                  {(reg58[(5'h13):(4'he)] || reg82[(4'h8):(2'h3)]),
                      (-(8'hbe))} : reg64) ~^ (wire32 || (~|(reg40[(3'h4):(3'h4)] ?
                  reg63[(3'h5):(3'h5)] : (reg77 ? reg54 : (8'hbc))))));
              reg82 <= ($signed($signed(reg82)) ?
                  reg24[(3'h4):(3'h4)] : $signed($signed({$unsigned(reg29),
                      (~&reg55)})));
              reg83 <= $unsigned($signed({(+$unsigned((8'hbb)))}));
              reg84 <= (|({$unsigned($signed(wire14))} || reg25[(3'h6):(3'h6)]));
            end
        end
    end
endmodule